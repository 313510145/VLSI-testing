
module dff (CK,RST,Q,D) ;
    input CK,RST,D ;
    output Q ;
    reg Q;
    always@(posedge CK)
    begin
	if(RST)
	    Q <= 1'd0 ;
	else
	    Q <= D ;
    end
endmodule

module s38584_seq(GND,VDD,CK,RST,g35,g36,g6744,g6745,g6746,g6747,g6748,g6749,g6750,
  g6751,g6752,g6753,g7243,g7245,g7257,g7260,g7540,g7916,g7946,g8132,g8178,g8215,g8235,
  g8277,g8279,g8283,g8291,g8342,g8344,g8353,g8358,g8398,g8403,g8416,g8475,g8719,g8783,
  g8784,g8785,g8786,g8787,g8788,g8789,g8839,g8870,g8915,g8916,g8917,g8918,g8919,g8920,
  g9019,g9048,g9251,g9497,g9553,g9555,g9615,g9617,g9680,g9682,g9741,g9743,g9817,g10122,
  g10306,g10500,g10527,g11349,g11388,g11418,g11447,g11678,g11770,g12184,g12238,g12300,
  g12350,g12368,g12422,g12470,g12832,g12919,g12923,g13039,g13049,g13068,g13085,g13099,
  g13259,g13272,g13865,g13881,g13895,g13906,g13926,g13966,g14096,g14125,g14147,g14167,
  g14189,g14201,g14217,g14421,g14451,g14518,g14597,g14635,g14662,g14673,g14694,g14705,
  g14738,g14749,g14779,g14828,g16603,g16624,g16627,g16656,g16659,g16686,g16693,g16718,
  g16722,g16744,g16748,g16775,g16874,g16924,g16955,g17291,g17316,g17320,g17400,g17404,
  g17423,g17519,g17577,g17580,g17604,g17607,g17639,g17646,g17649,g17674,g17678,g17685,
  g17688,g17711,g17715,g17722,g17739,g17743,g17760,g17764,g17778,g17787,g17813,g17819,
  g17845,g17871,g18092,g18094,g18095,g18096,g18097,g18098,g18099,g18100,g18101,g18881,
  g19334,g19357,g20049,g20557,g20652,g20654,g20763,g20899,g20901,g21176,g21245,g21270,
  g21292,g21698,g21727,g23002,g23190,g23612,g23652,g23683,g23759,g24151,g25114,g25167,
  g25219,g25259,g25582,g25583,g25584,g25585,g25586,g25587,g25588,g25589,g25590,g26801,
  g26875,g26876,g26877,g27831,g28030,g28041,g28042,g28753,g29210,g29211,g29212,g29213,
  g29214,g29215,g29216,g29217,g29218,g29219,g29220,g29221,g30327,g30329,g30330,g30331,
  g30332,g31521,g31656,g31665,g31793,g31860,g31861,g31862,g31863,g32185,g32429,g32454,
  g32975,g33079,g33435,g33533,g33636,g33659,g33874,g33894,g33935,g33945,g33946,g33947,
  g33948,g33949,g33950,g33959,g34201,g34221,g34232,g34233,g34234,g34235,g34236,g34237,
  g34238,g34239,g34240,g34383,g34425,g34435,g34436,g34437,g34597,g34788,g34839,g34913,
  g34915,g34917,g34919,g34921,g34923,g34925,g34927,g34956,g34972);
input GND,VDD,CK,RST,g35,g36,g6744,g6745,g6746,g6747,g6748,g6749,g6750,g6751,g6752,g6753;
output g7243,g7245,g7257,g7260,g7540,g7916,g7946,g8132,g8178,g8215,g8235,g8277,g8279,
  g8283,g8291,g8342,g8344,g8353,g8358,g8398,g8403,g8416,g8475,g8719,g8783,g8784,g8785,
  g8786,g8787,g8788,g8789,g8839,g8870,g8915,g8916,g8917,g8918,g8919,g8920,g9019,g9048,
  g9251,g9497,g9553,g9555,g9615,g9617,g9680,g9682,g9741,g9743,g9817,g10122,g10306,g10500,
  g10527,g11349,g11388,g11418,g11447,g11678,g11770,g12184,g12238,g12300,g12350,g12368,
  g12422,g12470,g12832,g12919,g12923,g13039,g13049,g13068,g13085,g13099,g13259,g13272,
  g13865,g13881,g13895,g13906,g13926,g13966,g14096,g14125,g14147,g14167,g14189,g14201,
  g14217,g14421,g14451,g14518,g14597,g14635,g14662,g14673,g14694,g14705,g14738,g14749,
  g14779,g14828,g16603,g16624,g16627,g16656,g16659,g16686,g16693,g16718,g16722,g16744,
  g16748,g16775,g16874,g16924,g16955,g17291,g17316,g17320,g17400,g17404,g17423,g17519,
  g17577,g17580,g17604,g17607,g17639,g17646,g17649,g17674,g17678,g17685,g17688,g17711,
  g17715,g17722,g17739,g17743,g17760,g17764,g17778,g17787,g17813,g17819,g17845,g17871,
  g18092,g18094,g18095,g18096,g18097,g18098,g18099,g18100,g18101,g18881,g19334,g19357,
  g20049,g20557,g20652,g20654,g20763,g20899,g20901,g21176,g21245,g21270,g21292,g21698,
  g21727,g23002,g23190,g23612,g23652,g23683,g23759,g24151,g25114,g25167,g25219,g25259,
  g25582,g25583,g25584,g25585,g25586,g25587,g25588,g25589,g25590,g26801,g26875,g26876,
  g26877,g27831,g28030,g28041,g28042,g28753,g29210,g29211,g29212,g29213,g29214,g29215,
  g29216,g29217,g29218,g29219,g29220,g29221,g30327,g30329,g30330,g30331,g30332,g31521,
  g31656,g31665,g31793,g31860,g31861,g31862,g31863,g32185,g32429,g32454,g32975,g33079,
  g33435,g33533,g33636,g33659,g33874,g33894,g33935,g33945,g33946,g33947,g33948,g33949,
  g33950,g33959,g34201,g34221,g34232,g34233,g34234,g34235,g34236,g34237,g34238,g34239,
  g34240,g34383,g34425,g34435,g34436,g34437,g34597,g34788,g34839,g34913,g34915,g34917,
  g34919,g34921,g34923,g34925,g34927,g34956,g34972;
  wire g72,g73,g84,g90,g91,g92,g99,g100,g110,g112,g113,g114,g115,g116,g120,g124,g125,g126,
    g127,g134,g135,g44,g45,g46,g47,g48,g49,g50,g51,g52,g53,g54,g55,g56,g57,g58,g63,g71,g85,g93,
    g101,g111,g43,g64,g65,g70,g4507,g4459,g4369,g4473,g4462,g4581,g4467,g4474,g4477,g4480,
    g4495,g4498,g4501,g4504,g4512,g4521,g4527,g4515,g4519,g4520,g4483,g4486,g4489,g4492,
    g4537,g4423,g4540,g4543,g4567,g4546,g4549,g4552,g4570,g4571,g4555,g4558,g4561,g4564,
    g4534,g4420,g4438,g4449,g4443,g4446,g4452,g4434,g4430,g4427,g4375,g4414,g4411,g4408,
    g4405,g4401,g4388,g4382,g4417,g4392,g4456,g4455,g1,g4304,g4308,g2932,g4639,g4621,g4628,
    g4633,g4643,g4340,g4349,g4358,g66,g4531,g4311,g4322,g4332,g4584,g4593,g4601,g4608,g4616,
    g4366,g4372,g4836,g4864,g4871,g4878,g4843,g4849,g4854,g4859,g4917,g4922,g4907,g4912,
    g4927,g4931,g4932,g4572,g4578,g4999,g5002,g5005,g5008,g4983,g4991,g4966,g4975,g4899,
    g4894,g4888,g4939,g4933,g4950,g4944,g4961,g4955,g4646,g4674,g4681,g4688,g4653,g4659,
    g4664,g4669,g4727,g4732,g4717,g4722,g4737,g4741,g4742,g59,g4575,g4809,g4812,g4815,g4818,
    g4793,g4801,g4776,g4785,g4709,g4704,g4698,g4749,g4743,g4760,g4754,g4771,g4765,g5313,
    g5290,g5320,g5276,g5283,g5308,g5327,g5331,g5335,g5339,g5343,g5348,g5352,g5357,g5297,
    g5101,g5109,g5062,g5105,g5112,g5022,g5016,g5029,g5033,g5037,g5041,g5046,g5052,g5057,
    g5069,g5073,g5077,g5080,g5084,g5092,g5097,g86,g5164,g5170,g5176,g5180,g5188,g5196,g5224,
    g5240,g5256,g5204,g5200,g5228,g5244,g5260,g5212,g5208,g5232,g5248,g5264,g5220,g5216,
    g5236,g5252,g5268,g5272,g128,g5156,g5120,g5115,g5124,g5128,g5134,g5138,g5142,g5148,
    g5152,g5160,g5659,g5637,g5666,g5623,g5630,g5654,g5673,g5677,g5681,g5685,g5689,g5694,
    g5698,g5703,g5644,g5448,g5456,g5406,g5452,g5459,g5366,g5360,g5373,g5377,g5381,g5385,
    g5390,g5396,g5401,g5413,g5417,g5421,g5424,g5428,g5436,g5441,g5445,g5511,g5517,g5523,
    g5527,g5535,g5543,g5571,g5587,g5603,g5551,g5547,g5575,g5591,g5607,g5559,g5555,g5579,
    g5595,g5611,g5567,g5563,g5583,g5599,g5615,g5619,g4821,g5503,g5467,g5462,g5471,g5475,
    g5481,g5485,g5489,g5495,g5499,g5507,g6005,g5983,g6012,g5969,g5976,g6000,g6019,g6023,
    g6027,g6031,g6035,g6040,g6044,g6049,g5990,g5794,g5802,g5752,g5798,g5805,g5712,g5706,
    g5719,g5723,g5727,g5731,g5736,g5742,g5747,g5759,g5763,g5767,g5770,g5774,g5782,g5787,
    g5791,g5857,g5863,g5869,g5873,g5881,g5889,g5917,g5933,g5949,g5897,g5893,g5921,g5937,
    g5953,g5905,g5901,g5925,g5941,g5957,g5913,g5909,g5929,g5945,g5961,g5965,g4831,g5849,
    g5813,g5808,g5817,g5821,g5827,g5831,g5835,g5841,g5845,g5853,g6351,g6329,g6358,g6315,
    g6322,g6346,g6365,g6369,g6373,g6377,g6381,g6386,g6390,g6395,g6336,g6140,g6148,g6098,
    g6144,g6151,g6058,g6052,g6065,g6069,g6073,g6077,g6082,g6088,g6093,g6105,g6109,g6113,
    g6116,g6120,g6128,g6133,g6137,g6203,g6209,g6215,g6219,g6227,g6235,g6263,g6279,g6295,
    g6243,g6239,g6267,g6283,g6299,g6251,g6247,g6271,g6287,g6303,g6259,g6255,g6275,g6291,
    g6307,g6311,g4826,g6195,g6159,g6154,g6163,g6167,g6173,g6177,g6181,g6187,g6191,g6199,
    g6697,g6675,g6704,g6661,g6668,g6692,g6711,g6715,g6719,g6723,g6727,g6732,g6736,g6741,
    g6682,g6486,g6494,g6444,g6490,g6497,g6404,g6398,g6411,g6415,g6419,g6423,g6428,g6434,
    g6439,g6451,g6455,g6459,g6462,g6466,g6474,g6479,g6483,g6549,g6555,g6561,g6565,g6573,
    g6581,g6609,g6625,g6641,g6589,g6585,g6613,g6629,g6645,g6597,g6593,g6617,g6633,g6649,
    g6605,g6601,g6621,g6637,g6653,g6657,g5011,g6541,g6505,g6500,g6509,g6513,g6519,g6523,
    g6527,g6533,g6537,g6545,g3303,g3281,g3310,g3267,g3274,g3298,g3317,g3321,g3325,g3329,
    g3338,g3343,g3347,g3352,g3288,g3092,g3100,g3050,g3096,g3103,g3010,g3004,g3017,g3021,
    g3025,g3029,g3034,g3040,g3045,g3057,g3061,g3065,g3068,g3072,g3080,g3085,g3089,g3155,
    g3161,g3167,g3171,g3179,g3187,g3215,g3231,g3247,g3195,g3191,g3219,g3235,g3251,g3203,
    g3199,g3223,g3239,g3255,g3211,g3207,g3227,g3243,g3259,g3263,g3333,g3147,g3111,g3106,
    g3115,g3119,g3125,g3129,g3133,g3139,g3143,g3151,g3654,g3632,g3661,g3618,g3625,g3649,
    g3668,g3672,g3676,g3680,g3689,g3694,g3698,g3703,g3639,g3443,g3451,g3401,g3447,g3454,
    g3361,g3355,g3368,g3372,g3376,g3380,g3385,g3391,g3396,g3408,g3412,g3416,g3419,g3423,
    g3431,g3436,g3440,g3506,g3512,g3518,g3522,g3530,g3538,g3566,g3582,g3598,g3546,g3542,
    g3570,g3586,g3602,g3554,g3550,g3574,g3590,g3606,g3562,g3558,g3578,g3594,g3610,g3614,
    g3684,g3498,g3462,g3457,g3466,g3470,g3476,g3480,g3484,g3490,g3494,g3502,g4005,g3983,
    g4012,g3969,g3976,g4000,g4019,g4023,g4027,g4031,g4040,g4045,g4049,g4054,g3990,g3794,
    g3802,g3752,g3798,g3805,g3712,g3706,g3719,g3723,g3727,g3731,g3736,g3742,g3747,g3759,
    g3763,g3767,g3770,g3774,g3782,g3787,g3791,g3857,g3863,g3869,g3873,g3881,g3889,g3917,
    g3933,g3949,g3897,g3893,g3921,g3937,g3953,g3905,g3901,g3925,g3941,g3957,g3913,g3909,
    g3929,g3945,g3961,g3965,g4035,g3849,g3813,g3808,g3817,g3821,g3827,g3831,g3835,g3841,
    g3845,g3853,g4165,g4169,g4125,g4072,g4064,g4057,g4141,g4082,g4076,g4087,g4093,g4098,
    g4108,g4104,g4145,g4112,g4116,g4119,g4122,g4153,g4164,g4129,g4132,g4135,g4138,g4172,
    g4176,g4146,g4157,g4258,g4264,g4269,g4273,g4239,g4294,g4297,g4300,g4253,g4249,g4245,
    g4277,g4281,g4284,g4287,g4291,g2946,g4191,g4188,g4194,g4197,g4200,g4204,g4207,g4210,
    g4180,g4185,g4213,g4216,g4219,g4222,g4226,g4229,g4232,g4235,g4242,g305,g311,g336,g324,
    g316,g319,g329,g333,g344,g347,g351,g355,g74,g106,g341,g637,g640,g559,g562,g568,g572,g586,
    g577,g582,g590,g595,g599,g604,g608,g613,g617,g622,g626,g632,g859,g869,g875,g878,g881,g884,
    g887,g872,g225,g255,g232,g262,g239,g269,g246,g446,g890,g862,g896,g901,g391,g365,g358,g370,
    g376,g385,g203,g854,g847,g703,g837,g843,g812,g817,g832,g822,g827,g723,g645,g681,g699,g650,
    g655,g718,g661,g728,g79,g691,g686,g667,g671,g676,g714,g499,g504,g513,g518,g528,g482,g490,
    g417,g411,g424,g475,g441,g437,g433,g429,g401,g392,g405,g182,g174,g168,g460,g452,g457,g471,
    g464,g468,g479,g102,g496,g732,g753,g799,g802,g736,g739,g744,g749,g758,g763,g767,g772,g776,
    g781,g785,g790,g794,g807,g554,g538,g546,g542,g534,g550,g136,g199,g278,g283,g287,g291,g294,
    g298,g142,g146,g164,g150,g153,g157,g160,g301,g222,g194,g191,g209,g215,g218,g1249,g1266,
    g1280,g1252,g1256,g1259,g1263,g1270,g1274,g1277,g1418,g1422,g1426,g1430,g1548,g1564,
    g1559,g1554,g1570,g1585,g1589,g1576,g1579,g1339,g1500,g1582,g1333,g1399,g1459,g1322,
    g1514,g1526,g1521,g1306,g1532,g1536,g1542,g1413,g1395,g1404,g1319,g1312,g1351,g1345,
    g1361,g1367,g1373,g1379,g1384,g1389,g1489,g1495,g1442,g1437,g1478,g1454,g1448,g1467,
    g1472,g1484,g1300,g1291,g1296,g1283,g1287,g1311,g929,g904,g921,g936,g907,g911,g914,g918,
    g925,g930,g933,g1075,g1079,g1083,g1087,g1205,g1221,g1216,g1211,g1227,g1242,g1246,g1233,
    g1236,g996,g1157,g1239,g990,g1056,g1116,g979,g1171,g1183,g1178,g962,g1189,g1193,g1199,
    g1070,g1052,g1061,g976,g969,g1008,g1002,g1018,g1024,g1030,g1036,g1041,g1046,g1146,g1152,
    g1099,g1094,g1135,g1111,g1105,g1124,g1129,g1141,g956,g947,g952,g939,g943,g967,g968,g1592,
    g1644,g1636,g1668,g1682,g1687,g1604,g1600,g1608,g1620,g1616,g1612,g1632,g1624,g1648,
    g1664,g1657,g1677,g1691,g1696,g1700,g1706,g1710,g1714,g1720,g1724,g1728,g1779,g1772,
    g1802,g1816,g1821,g1740,g1736,g1744,g1756,g1752,g1748,g1768,g1760,g1783,g1798,g1792,
    g1811,g1825,g1830,g1834,g1840,g1844,g1848,g1854,g1858,g1862,g1913,g1906,g1936,g1950,
    g1955,g1874,g1870,g1878,g1890,g1886,g1882,g1902,g1894,g1917,g1932,g1926,g1945,g1959,
    g1964,g1968,g1974,g1978,g1982,g1988,g1992,g1996,g2047,g2040,g2070,g2084,g2089,g2008,
    g2004,g2012,g2024,g2020,g2016,g2036,g2028,g2051,g2066,g2060,g2079,g2093,g2098,g2102,
    g2108,g2112,g2116,g2122,g2126,g2130,g2138,g2145,g2151,g2152,g2153,g2204,g2197,g2227,
    g2241,g2246,g2165,g2161,g2169,g2181,g2177,g2173,g2193,g2185,g2208,g2223,g2217,g2236,
    g2250,g2255,g2259,g2265,g2269,g2273,g2279,g2283,g2287,g2338,g2331,g2361,g2375,g2380,
    g2299,g2295,g2303,g2315,g2311,g2307,g2327,g2319,g2342,g2357,g2351,g2370,g2384,g2389,
    g2393,g2399,g2403,g2407,g2413,g2417,g2421,g2472,g2465,g2495,g2509,g2514,g2433,g2429,
    g2437,g2449,g2445,g2441,g2461,g2453,g2476,g2491,g2485,g2504,g2518,g2523,g2527,g2533,
    g2537,g2541,g2547,g2551,g2555,g2606,g2599,g2629,g2643,g2648,g2567,g2563,g2571,g2583,
    g2579,g2575,g2595,g2587,g2610,g2625,g2619,g2638,g2652,g2657,g2661,g2667,g2671,g2675,
    g2681,g2685,g2689,g2697,g2704,g2710,g2711,g2837,g2841,g2712,g2715,g2719,g2724,g2729,
    g2735,g2741,g2748,g2756,g2759,g2763,g2767,g2779,g2791,g2795,g2787,g2783,g2775,g2771,
    g2831,g121,g2799,g2811,g2823,g2827,g2819,g2815,g2807,g2803,g2834,g117,g2999,g2994,g2988,
    g2868,g2873,g2890,g2844,g2852,g2860,g2894,g37,g94,g2848,g2856,g2864,g2898,g2882,g2878,
    g2886,g2980,g2984,g2907,g2912,g2922,g2936,g2950,g2960,g2970,g2902,g2917,g2927,g2941,
    g2955,g2965,g2975,g3003,g5,g6,g7,g8,g9,g16,g19,g28,g31,g34,g12,g22,g25,I11617,g6754,I11620,
    g6755,I11623,g6756,I11626,g6767,I11629,g6772,I11632,g6782,I11635,g6789,g6799,g6800,
    g6801,g6802,g6803,g6804,g6808,g6809,g6810,g6811,g6814,g6815,g6816,g6817,g6818,g6819,
    g6820,I11655,g6821,g6825,g6826,g6827,g6828,g6829,g6830,g6831,I11665,g6832,g6836,g6837,
    g6838,g6839,g6840,g6841,g6845,g6846,g6847,g6848,g6849,g6850,g6854,g6855,I11682,g6856,
    I11685,g6867,I11688,g6868,I11691,g6869,g6870,g6873,g6874,I11697,g6875,g6887,I11701,
    g6888,g6895,g6900,g6903,g6904,I11708,g6905,g6917,g6918,g6923,g6926,g6927,I11716,g6928,
    g6940,g6941,I11721,g6946,g6953,g6954,I11726,g6955,g6956,g6957,g6958,g6959,g6960,I11734,
    g6961,I11737,g6971,I11740,g6972,I11743,g6973,I11746,g6974,g6975,I11750,g6976,I11753,
    g6977,g6978,g6982,g6983,g6984,g6985,g6986,g6987,g6988,g6989,g6990,g6991,g6992,g6993,
    g6994,g6995,g6996,g6997,g6998,g6999,g7002,g7003,I11777,g7004,g7017,g7018,g7023,g7026,
    g7027,I11785,g7028,g7040,g7041,g7046,g7049,g7050,I11793,g7051,g7063,g7064,g7069,g7072,
    g7073,I11801,g7074,g7086,g7087,g7092,g7095,g7096,I11809,g7097,g7109,g7110,g7115,g7116,
    I11816,g7117,g7118,I11820,g7121,g7132,g7134,g7138,I11835,g7148,g7149,g7153,g7157,I11843,
    g7161,g7162,g7163,g7166,g7170,g7174,g7178,g7183,g7187,g7191,g7195,I11860,g7196,g7197,
    g7202,g7212,g7216,g7219,g7222,g7224,g7231,g7232,g7235,g7236,g7239,I11892,g7244,I11896,
    g7246,g7247,g7252,I11903,g7258,g7259,I11908,g7261,g7262,g7266,g7267,g7268,g7275,g7280,
    g7285,g7289,g7293,g7296,g7297,g7301,g7308,g7314,g7315,g7322,g7327,g7328,g7335,g7340,
    g7343,g7344,g7345,g7349,g7356,g7361,g7362,g7369,g7374,g7379,g7380,g7387,g7392,g7393,
    g7394,g7395,g7397,g7400,g7405,g7410,g7411,g7418,g7423,g7424,g7431,g7436,g7437,g7438,
    g7439,g7440,g7441,g7443,g7446,g7451,g7456,g7461,g7462,g7470,g7471,g7472,g7473,I11980,
    g7474,g7475,g7479,g7487,g7490,g7495,g7496,g7497,g7498,I11992,g7502,g7503,g7512,g7513,
    g7514,I12000,g7515,I12003,g7516,g7517,g7518,g7519,g7521,g7522,g7523,I12013,g7526,
    I12016,g7527,g7528,g7532,g7533,g7534,g7535,g7536,g7537,I12026,g7541,I12030,g7542,I12033,
    g7543,g7544,g7548,g7553,g7557,I12041,g7558,g7563,g7564,I12046,g7565,I12049,g7566,g7577,
    g7581,I12056,g7586,g7591,g7592,I12061,g7593,I12064,g7594,I12067,g7595,I12070,g7596,
    g7597,I12083,g7615,I12086,g7616,I12089,g7617,I12092,g7618,g7619,I12103,g7623,I12106,
    g7624,I12109,g7625,I12112,g7626,g7627,g7631,I12117,g7632,I12120,g7633,I12123,g7634,
    g7635,g7636,I12128,g7640,g7643,I12132,g7647,I12135,g7648,g7649,g7650,g7655,I12141,
    g7659,I12144,g7660,g7666,g7670,I12151,g7674,g7680,g7686,I12159,g7689,g7693,g7697,
    I12167,g7704,g7715,g7716,I12172,g7717,g7733,I12176,g7738,g7749,g7750,g7751,g7752,I12183,
    g7753,g7765,I12189,g7766,g7778,g7779,g7780,g7785,g7788,I12199,g7791,g7802,g7805,g7806,
    g7809,I12214,g7812,g7824,g7827,g7828,I12227,g7831,g7835,g7840,g7841,g7845,g7851,g7854,
    g7858,g7863,g7867,g7868,g7870,g7873,g7876,g7880,g7886,g7888,g7891,g7892,g7898,g7903,
    g7907,g7908,g7909,g7913,I12300,g7917,g7922,g7926,g7927,g7928,g7933,g7936,g7939,g7943,
    I12314,g7947,g7952,g7953,g7957,g7960,g7963,g7964,g7970,g7971,g7972,g7975,g7980,g7985,
    g7991,g7992,I12333,g7993,I12336,g7994,g7995,g7998,g8002,g8005,g8009,g8011,g8016,g8021,
    g8026,I12355,g8032,g8033,g8037,I12360,g8038,g8046,g8052,g8055,g8056,g8057,g8058,g8059,
    g8064,g8068,g8070,g8075,g8080,I12382,g8085,g8087,g8088,g8091,g8092,g8093,g8097,g8102,
    g8106,g8107,g8112,g8113,g8114,g8119,g8123,g8125,g8130,I12411,g8133,I12415,g8134,I12418,
    g8135,g8136,g8137,g8138,g8139,g8146,g8150,g8154,g8155,g8160,g8164,g8165,g8170,g8171,
    g8172,I12437,g8179,g8180,g8181,g8183,g8186,g8187,g8195,g8201,g8205,g8211,I12451,g8216,
    g8217,g8218,g8219,g8224,g8228,g8229,I12463,g8236,g8237,g8239,g8240,g8241,g8249,g8255,
    g8259,g8267,g8273,I12483,g8278,I12487,g8280,g8281,g8282,I12493,g8284,I12497,g8285,
    g8286,g8287,g8290,I12503,g8296,g8297,g8300,g8301,g8302,g8310,g8316,g8324,g8330,g8334,
    g8340,g8341,I12519,g8343,I12523,g8345,g8346,g8350,I12530,g8354,I12534,g8355,g8356,
    I12538,g8357,I12541,g8362,g8363,g8364,g8365,g8373,g8381,g8387,g8388,g8389,g8390,g8396,
    g8397,I12563,g8399,g8400,I12568,g8404,I12572,g8405,g8406,g8407,I12577,g8411,I12580,
    g8418,g8426,g8431,g8438,g8439,g8440,g8441,g8442,g8443,g8449,g8450,g8451,g8456,g8457,
    g8458,g8462,g8466,I12605,g8470,I12608,g8477,g8478,g8479,g8480,I12618,g8481,g8492,g8497,
    g8504,g8505,g8506,g8507,g8508,g8509,g8514,I12631,g8515,g8519,g8522,g8526,g8531,g8534,
    g8538,g8539,g8540,g8541,I12644,g8542,g8553,g8558,g8565,g8566,g8567,g8571,I12654,g8572,
    g8575,g8579,g8584,g8587,g8591,g8592,g8593,g8594,I12666,g8595,g8606,g8607,g8608,g8612,
    g8616,g8620,g8623,g8626,g8630,g8631,g8635,g8639,g8644,g8647,g8650,g8651,g8654,g8655,
    g8659,g8663,g8666,g8669,g8672,g8673,g8676,g8677,g8680,g8681,g8685,g8686,g8696,g8697,
    g8700,I12709,g8703,I12712,g8712,g8713,g8714,g8715,g8718,I12719,g8725,g8733,g8734,
    I12735,g8740,g8741,g8742,g8743,g8744,g8745,g8748,g8756,I12746,g8757,I12749,g8763,g8764,
    g8765,g8766,g8770,g8774,I12758,g8778,I12761,I12764,I12767,I12770,I12773,I12776,I12779,
    I12787,g8791,I12790,g8792,I12793,g8795,g8796,g8804,I12799,g8805,g8807,g8808,I12805,
    g8812,I12808,g8818,I12811,g8821,g8822,g8830,g8833,g8836,I12819,g8840,I12823,g8841,
    I12826,g8844,g8848,g8851,g8854,g8858,g8859,I12837,g8872,I12855,g8876,I12858,g8879,
    I12861,g8880,g8883,g8890,g8891,g8895,g8898,g8899,g8903,g8912,g8914,I12884,I12887,I12890,
    I12893,I12896,I12899,I12907,g8922,I12910,g8925,g8928,g8938,g8944,g8945,g8948,g8951,
    g8954,g8955,g8964,I12927,g8971,I12930,g8974,g8977,I12935,g8989,g8990,g8993,g8997,g9000,
    g9003,g9007,g9011,g9014,g9018,I12950,g9020,I12954,g9021,g9024,g9030,g9036,g9037,g9040,
    g9044,I12963,g9049,g9050,g9051,g9056,g9060,g9064,g9070,g9071,g9072,g9073,g9077,g9083,
    g9086,g9091,g9095,g9099,g9103,I12987,g9104,g9152,I12991,g9153,I12994,g9154,I12997,
    g9155,g9158,g9162,g9166,g9174,g9180,g9184,I13007,g9185,I13010,g9186,g9187,g9194,g9197,
    g9200,g9206,g9212,I13020,g9213,g9214,g9220,g9223,g9226,g9229,g9234,g9239,I13031,g9245,
    g9247,g9250,I13037,g9252,g9253,g9257,g9259,g9264,g9269,g9274,I13054,g9280,I13057,g9281,
    g9282,g9283,g9284,g9285,g9291,g9298,g9299,g9300,g9305,g9309,g9311,g9316,g9321,g9326,
    g9332,g9333,g9337,g9338,g9339,I13094,g9340,g9354,g9360,g9364,g9369,g9373,g9374,g9379,
    g9380,g9381,g9386,g9390,g9392,g9397,g9402,g9407,g9413,g9414,g9415,g9416,I13124,g9417,
    g9429,g9433,g9434,g9439,g9443,g9444,g9449,g9450,g9451,g9456,g9460,g9462,g9467,g9472,
    I13149,g9477,I13152,g9478,g9480,g9484,g9488,g9489,g9490,g9491,g9492,g9496,I13166,g9498,
    g9499,g9500,g9501,g9506,g9510,g9511,g9516,g9517,g9518,g9523,g9527,g9529,g9534,g9537,
    g9541,g9542,g9546,g9547,g9551,g9552,I13202,g9554,I13206,g9556,g9557,g9558,g9559,g9564,
    g9568,g9569,g9574,g9575,g9576,g9581,g9582,g9585,g9590,g9594,g9598,g9599,g9600,g9601,
    g9607,g9613,g9614,I13236,g9616,I13240,g9618,g9619,g9620,g9621,g9626,g9630,g9631,g9636,
    I13252,g9637,g9638,g9639,g9644,g9648,g9653,g9657,g9660,g9661,g9662,g9669,g9670,g9671,
    g9672,g9678,g9679,I13276,g9681,I13280,g9683,g9684,g9685,g9686,I13287,g9687,g9688,g9689,
    g9690,g9691,g9692,g9693,g9698,g9699,g9704,g9708,g9713,g9714,g9716,g9721,g9728,g9729,
    g9730,g9731,g9732,g9733,g9739,g9740,I13317,g9742,I13321,g9744,g9745,I13326,g9746,
    I13329,g9747,g9748,g9749,g9751,g9752,g9753,g9754,g9759,g9760,g9761,g9766,g9771,I13352,
    g9772,g9776,g9777,g9778,g9779,I13360,g9780,g9792,g9797,g9804,g9805,g9806,g9807,g9808,
    g9809,g9815,g9816,I13374,g9818,g9819,g9820,g9821,g9822,g9824,g9826,g9827,g9828,g9829,
    g9831,g9832,g9833,g9834,g9839,g9842,g9843,g9848,g9853,g9856,g9860,g9861,g9862,g9863,
    I13424,g9864,g9875,g9880,g9887,g9888,g9889,g9890,g9891,g9892,g9898,g9899,g9900,g9901,
    g9902,g9903,g9905,g9907,g9909,g9910,g9911,g9913,g9914,g9915,g9916,I13473,g9917,g9920,
    g9924,g9927,g9931,g9932,g9933,g9934,I13483,g9935,g9946,g9951,g9958,g9959,g9960,g9961,
    g9962,g9963,g9964,g9965,g9969,g9970,g9971,g9973,g9974,g9976,g9977,g9978,g9982,g9983,
    g9985,g9989,g9992,g9995,g9999,g10000,g10001,g10002,I13539,g10003,g10014,g10019,g10026,
    g10027,g10028,I13548,g10029,g10030,I13552,g10031,g10032,g10033,g10035,g10036,g10037,
    g10038,g10039,g10040,g10042,g10043,g10044,g10047,g10050,g10053,g10057,g10058,g10059,
    g10060,I13581,g10061,g10072,g10073,g10074,g10077,g10078,g10079,g10080,g10081,g10082,
    g10083,g10084,g10085,g10086,I13597,g10087,g10090,g10093,g10096,g10099,g10102,g10106,
    I13606,g10107,g10108,g10109,g10110,g10111,g10112,g10113,g10114,g10115,g10116,g10117,
    g10118,g10119,g10120,g10121,I13623,g10129,g10130,g10133,g10136,g10139,g10140,I13634,
    g10141,I13637,g10142,g10143,g10147,g10150,g10151,g10152,g10153,g10154,g10155,g10156,
    g10157,g10158,g10159,g10165,g10166,g10169,g10172,g10175,g10176,g10177,g10178,g10180,
    g10181,g10182,g10183,g10184,g10190,g10191,g10194,g10197,I13672,g10198,g10199,g10200,
    g10203,g10204,g10206,g10212,g10213,I13684,g10216,g10217,g10218,g10219,g10222,g10223,
    g10229,I13694,g10230,g10231,g10232,I13699,g10233,g10261,g10262,I13705,g10272,I13708,
    g10273,g10274,g10275,g10278,I13715,g10287,I13718,g10288,g10289,I13723,g10295,I13726,
    g10308,g10311,I13740,g10319,g10320,I13744,g10323,g10334,g10335,g10337,I13759,g10347,
    I13762,g10348,g10349,g10350,g10351,g10352,g10353,g10354,g10355,g10356,g10357,g10358,
    g10359,g10360,g10361,g10362,I13779,g10363,g10364,g10365,g10366,g10367,g10368,g10369,
    g10370,g10371,g10372,g10373,g10374,g10375,g10376,g10377,g10378,g10379,g10380,g10381,
    g10382,g10383,I13802,g10384,I13805,g10385,g10386,g10387,g10388,g10389,g10390,g10391,
    g10392,g10393,g10394,g10395,g10396,g10397,g10398,g10399,g10400,g10401,g10402,g10403,
    g10404,g10405,g10406,g10407,g10408,g10409,g10410,g10411,g10412,g10413,g10414,g10415,
    g10416,g10417,g10418,g10419,g10420,g10427,g10428,g10429,I13847,g10430,I13857,g10473,
    g10474,g10475,g10487,g10489,g10490,g10497,g10498,I13872,g10499,I13875,g10502,g10503,
    g10504,g10509,g10518,g10519,I13889,g10521,I13892,g10530,g10531,g10532,g10533,g10540,
    g10541,g10542,I13906,g10544,g10553,g10554,g10564,g10570,g10571,g10572,g10581,g10582,
    g10597,g10606,g10607,g10608,g10612,g10613,g10620,g10621,I13968,g10627,g10652,I13979,
    g10658,g10664,I13990,g10678,I13995,g10685,g10708,I14006,g10710,g10725,I14016,g10727,
    g10741,g10761,g10762,I14033,g10776,g10794,g10795,g10804,I14046,g10805,I14050,g10812,
    g10815,I14054,g10816,g10830,I14069,g10851,g10857,g10872,I14079,g10877,g10881,g10882,
    g10897,g10960,g10980,I14119,g10981,g11011,g11017,g11026,g11030,g11031,g11033,g11034,
    g11038,g11042,g11043,I14158,g11048,g11110,g11122,g11128,g11129,I14192,g11136,g11143,
    g11147,g11164,I14222,g11165,g11170,g11181,I14241,g11182,g11183,g11192,I14267,g11202,
    I14271,g11204,g11214,g11215,g11233,g11234,I14301,g11235,g11236,I14305,g11237,g11249,
    g11250,g11268,g11269,I14326,g11290,g11291,g11293,g11294,g11316,I14346,g11317,g11324,
    g11325,g11336,g11344,I14365,I14381,g11367,g11371,g11373,g11383,I14395,I14409,g11398,
    g11401,g11402,g11403,g11404,g11413,I14424,g11425,g11428,g11429,g11430,g11431,I14450,
    I14455,g11450,g11467,g11468,g11470,g11471,g11472,I14475,g11498,g11509,g11510,g11512,
    g11513,g11519,I14505,g11547,g11560,g11562,g11576,I14537,g11592,g11608,g11609,g11615,
    g11631,I14550,g11640,g11652,g11663,g11677,I14563,I14567,g11686,I14570,g11691,g11702,
    I14576,g11705,I14579,g11706,I14584,g11709,g11714,I14589,g11720,g11721,I14593,g11724,
    g11735,g11736,g11741,I14602,g11744,g11753,g11754,g11762,g11769,I14619,I14623,g11772,
    g11779,g11786,I14630,g11790,I14633,g11793,g11796,g11810,g11811,g11812,g11815,g11819,
    I14644,g11820,I14647,g11823,I14650,g11826,I14653,g11829,g11832,g11833,g11841,I14660,
    g11842,I14663,g11845,g11849,I14668,g11852,I14671,g11855,g11861,g11865,g11866,I14679,
    g11867,g11868,I14684,g11872,I14687,g11875,I14690,g11878,g11884,g11888,g11889,I14702,
    g11894,I14705,g11897,I14708,g11900,g11910,g11911,g11912,I14727,g11917,I14730,g11920,
    g11927,I14742,g11928,I14745,g11929,g11930,I14749,g11931,I14761,g11941,g11948,I14773,
    g11949,g11963,g11964,I14797,g11965,I14800,g11966,I14823,g11981,g11984,I14827,g11985,
    I14830,g11986,I14833,g11987,I14836,g11988,I14839,g11989,g11991,I14862,g12009,g12012,
    I14866,g12013,g12018,g12021,g12036,I14893,g12037,I14896,g12038,I14899,g12039,I14902,
    g12040,I14905,g12041,g12047,g12051,g12054,I14932,g12074,I14935,g12075,g12076,I14939,
    g12077,g12082,g12086,g12088,g12107,I14964,g12108,I14967,g12109,I14970,g12110,g12122,
    I14999,g12143,g12180,g12181,I15030,g12182,I15033,g12183,I15036,I15070,g12217,I15073,
    g12218,g12233,I15102,g12295,I15144,g12321,I15162,g12322,g12337,g12345,I15190,I15205,
    g12367,I15208,g12378,I15223,g12381,g12399,g12417,I15238,I15250,g12430,g12440,g12465,
    I15284,I15295,g12477,g12487,I15316,g12490,g12497,g12543,g12546,g12563,g12598,g12614,
    I15382,g12640,g12656,g12672,g12705,g12721,g12738,g12749,g12760,g12778,g12779,g12790,
    g12793,g12804,g12805,g12811,g12818,g12820,g12823,g12830,g12831,I15448,g12833,g12834,
    g12835,g12836,g12837,g12838,g12839,g12840,g12841,g12842,g12843,g12844,g12845,I15474,
    g12857,g12859,g12860,g12861,g12862,g12863,g12864,g12865,g12866,g12867,g12868,g12869,
    g12870,g12871,g12872,g12873,g12874,I15494,g12875,g12878,g12879,g12880,g12881,g12882,
    g12883,g12884,g12885,g12886,g12887,g12888,g12889,g12890,g12891,g12892,g12893,g12894,
    g12895,g12896,g12897,g12898,g12899,g12900,g12901,g12902,g12903,g12904,g12905,g12906,
    g12907,g12908,g12909,g12914,I15533,g12918,I15536,g12921,g12922,I15542,g12929,g12930,
    I15550,g12932,g12936,g12937,I15556,g12938,g12940,g12944,g12945,I15564,g12946,g12950,
    I15569,g12951,I15572,g12952,I15577,g12955,g12967,g12968,g12975,I15587,g12976,I15590,
    g12977,I15593,g12978,I15600,g12983,g12995,g12996,g12997,g12998,I15609,g13003,g13007,
    g13008,I15617,g13009,I15620,g13010,I15623,g13011,I15626,g13012,g13014,g13015,g13016,
    I15633,g13017,I15636,g13018,g13022,g13023,g13024,g13026,I15647,g13027,I15650,g13028,
    g13033,g13034,g13036,g13037,I15663,I15667,g13041,g13045,I15677,g13051,I15682,g13055,
    g13061,g13062,g13064,g13065,I15697,g13070,I15702,g13074,I15705,g13075,g13082,I15717,
    g13087,I15727,g13096,I15732,I15736,g13101,g13103,g13106,g13107,g13116,g13117,g13120,
    g13132,g13133,I15765,g13138,g13140,g13141,g13142,I15773,g13144,g13173,g13174,g13175,
    I15782,g13177,g13188,g13189,g13190,I15788,g13191,g13209,g13215,g13216,g13222,I15800,
    g13223,g13239,g13246,g13249,I15811,g13250,I15814,g13251,g13255,I15821,g13258,I15824,
    I15831,g13267,I15834,g13271,I15837,g13278,I15843,g13279,I15846,g13280,g13297,I15862,
    g13298,g13301,g13302,I15869,g13303,I15872,g13304,g13305,I15878,g13311,g13312,g13314,
    g13322,g13323,I15893,g13329,g13334,I15906,g13350,I15915,g13394,I15918,g13409,I15921,
    g13410,g13412,g13413,g13414,I15929,g13416,I15932,g13431,I15937,g13437,g13458,I15942,
    g13460,g13463,g13474,I15954,g13477,g13483,g13484,g13485,g13494,g13504,g13505,g13506,
    I15981,g13510,I15987,g13514,g13521,g13522,g13530,I16010,g13545,g13555,g13565,g13569,
    I16024,g13574,I16028,g13583,g13584,g13593,g13594,g13595,g13596,I16040,g13605,g13620,
    g13621,g13624,g13625,g13626,g13637,I16057,g13638,g13655,g13663,g13664,g13665,g13675,
    g13679,I16077,g13680,g13706,g13707,g13715,I16090,g13716,g13729,g13736,I16102,g13745,
    g13763,I16117,g13782,I16120,g13793,I16135,g13809,I16150,g13835,I16160,g13856,I16163,
    g13857,I16168,g13868,g13869,g13876,g13877,I16181,g13885,I16193,g13901,g13902,I16201,
    I16217,g13932,g13933,I16231,g13943,I16246,g13975,g13976,g13995,g13999,g14004,g14029,
    I16289,g14031,g14032,g14034,g14063,g14065,g14095,I16328,I16345,I16357,g14149,g14150,
    g14166,I16371,g14169,g14173,g14179,g14183,g14184,g14186,I16391,g14191,g14192,g14197,
    g14198,I16401,g14203,g14204,g14205,g14208,g14209,g14215,I16417,g14219,g14226,g14231,
    g14232,g14237,g14238,g14251,I16438,g14252,g14255,g14262,g14275,I16452,g14276,I16455,
    g14277,I16460,g14290,g14297,I16468,g14307,I16471,g14308,I16476,g14314,I16479,g14315,
    g14321,I16486,g14330,I16489,g14331,I16492,g14332,I16498,g14336,I16502,g14338,g14342,
    g14348,g14357,I16512,g14358,I16515,g14359,I16521,g14363,I16526,g14366,g14376,g14377,
    I16535,g14383,I16538,g14384,I16541,g14385,I16544,g14386,I16555,g14398,g14405,g14406,
    I16564,g14412,I16575,I16579,g14423,g14424,g14431,g14432,I16590,g14441,I16593,g14442,
    I16596,g14443,I16606,I16610,g14453,I16613,g14454,g14503,g14504,I16626,g14509,I16629,
    g14510,I16639,g14535,I16651,g14536,g14541,I16660,g14543,I16663,g14544,g14545,g14562,
    I16676,g14563,I16679,g14564,I16688,g14571,I16698,g14582,g14584,I16709,g14591,I16713,
    I16724,g14609,I16733,g14616,g14630,g14631,I16741,I16747,g14639,I16755,g14645,I16762,
    g14668,g14669,I16770,I16775,g14676,I16795,g14700,g14701,I16803,g14714,I16821,g14744,
    g14745,I16829,g14753,I16847,g14785,g14786,I16855,g14790,I16875,g14833,I16898,g14873,
    I16917,g14912,I16969,g15048,I17008,g15085,I17094,g15169,I17098,g15171,I17101,g15224,
    I17104,g15277,g15344,I17108,g15345,I17111,g15348,I17114,g15371,I17118,g15373,I17121,
    g15426,g15479,I17125,g15480,I17128,g15483,I17131,g15506,I17136,g15509,g15562,I17140,
    g15563,I17143,g15566,g15568,I17148,g15569,g15571,I17154,g15573,I17159,g15579,g15580,
    I17166,g15588,I17173,g15595,g15614,I17181,g15615,I17188,g15634,g15655,I17198,g15656,
    I17207,g15680,g15705,I17228,g15714,g15731,I17249,g15733,g15739,g15740,g15746,g15747,
    g15750,g15755,g15756,I17276,g15758,g15799,I17302,g15806,g15811,I17314,g15816,I17324,
    g15824,g15830,g15831,g15842,I17355,g15862,I17374,g15885,I17392,g15915,I17395,g15932,
    I17401,g15938,I17416,g15969,I17420,g15979,I17425,g16000,g16030,I17436,g16031,I17442,
    g16053,g16075,I17456,g16077,g16096,g16099,I17471,g16100,g16123,g16124,g16127,I17488,
    g16129,I17491,g16136,g16158,g16159,g16162,I17507,g16164,g16171,g16172,g16180,g16182,
    g16186,g16195,g16197,g16200,g16206,g16214,I17557,g16216,g16223,I17569,g16228,g16235,
    I17590,g16249,g16280,I17609,g16284,I17612,g16285,I17615,g16286,g16289,g16290,I17626,
    g16300,g16305,I17633,g16307,I17636,g16308,I17639,g16309,g16310,g16311,g16320,I17650,
    g16322,I17653,g16323,g16325,I17658,g16326,I17661,g16349,g16423,I17668,g16428,I17671,
    g16429,I17675,g16431,I17679,g16449,g16472,g16473,g16475,g16482,I17695,g16487,I17699,
    g16489,I17704,g16508,g16509,g16510,g16511,g16512,g16514,g16515,g16521,g16522,g16523,
    I17723,g16525,g16526,g16527,g16528,g16529,g16530,I17733,g16533,I17744,g16540,I17747,
    g16577,I17750,g16578,g16579,I17754,g16580,g16582,g16583,g16584,g16585,I17763,g16587,
    g16588,g16589,I17772,g16594,I17780,g16600,I17783,g16601,g16602,I17787,g16605,g16606,
    g16607,g16608,g16609,I17801,g16615,I17808,g16620,g16622,g16623,I17814,g16626,I17819,
    g16629,g16630,g16631,g16632,I17834,g16640,I17839,g16643,I17842,g16644,g16645,g16651,
    g16652,g16654,g16655,I17852,g16658,I17857,g16661,I17873,g16675,I17876,g16676,I17879,
    g16677,g16680,g16684,g16685,I17892,g16688,g16689,g16691,g16692,I17901,g16695,I17916,
    g16708,I17919,g16709,g16712,g16716,g16717,I17932,g16720,g16721,I17938,g16724,g16725,
    g16726,g16727,I17956,g16738,g16739,g16740,g16742,g16743,I17964,g16746,g16747,I17970,
    g16750,I17976,g16752,I17989,g16767,g16768,g16769,g16771,g16773,g16774,I17999,I18003,
    g16777,I18006,g16782,I18009,g16795,g16809,g16812,g16814,I18028,g16816,I18031,g16821,
    I18034,g16826,g16853,I18048,g16856,I18051,g16861,I18060,g16872,I18063,g16873,I18066,
    I18071,g16877,I18078,g16886,I18083,g16897,I18086,g16920,I18089,g16923,I18092,I18101,
    g16931,I18104,g16954,I18107,g16958,I18114,g16960,I18117,g16963,I18120,g16964,g16966,
    I18125,g16967,g16968,g16969,I18131,g16971,I18135,g16987,I18138,g17010,g17013,g17014,
    I18143,g17015,g17056,I18148,g17058,I18151,g17059,I18154,g17062,g17085,g17086,g17087,
    I18160,g17088,g17092,I18165,g17093,I18168,g17096,g17120,g17121,g17122,g17124,I18177,
    g17125,I18180,g17128,g17135,g17136,I18191,g17141,g17144,g17147,g17154,I18205,g17155,
    g17157,I18214,g17178,I18221,g17183,I18224,g17188,g17189,I18233,g17197,I18238,g17200,
    g17216,I18245,g17221,I18248,g17224,I18252,g17226,g17242,I18259,g17247,I18262,g17248,
    I18265,g17249,I18270,g17271,I18276,I18280,g17296,g17301,I18285,g17302,g17308,I18293,
    I18297,I18301,g17324,I18304,g17325,I18307,g17326,I18310,g17327,I18313,g17328,g17366,
    I18320,g17367,I18323,g17384,g17389,g17390,g17392,I18333,I18337,I18341,g17408,I18344,
    g17409,g17410,g17411,I18350,g17413,g17414,g17415,g17416,g17417,g17419,I18360,I18364,
    g17427,I18367,g17428,I18370,g17429,I18373,g17430,I18376,g17431,I18379,g17432,I18382,
    g17433,g17465,g17466,g17467,g17470,g17471,g17472,g17473,I18398,g17475,g17476,g17477,
    g17478,g17479,g17481,I18408,g17485,I18411,g17486,I18414,g17487,g17489,g17491,g17494,
    g17496,g17497,g17498,g17499,I18434,g17501,g17502,g17503,g17504,g17505,g17507,I18443,
    g17508,I18446,g17509,g17512,g17518,I18460,g17521,g17522,g17523,g17524,I18469,g17526,
    g17527,g17528,g17529,g17530,I18476,g17531,I18479,g17532,I18482,g17533,g17573,g17575,
    g17576,I18504,g17579,I18509,g17582,g17583,g17584,g17585,I18518,g17587,g17588,g17589,
    I18523,g17590,I18526,g17591,g17599,g17600,g17602,g17603,I18555,g17606,I18560,g17609,
    g17610,g17611,g17612,I18571,g17614,I18574,g17615,g17616,g17637,g17638,I18600,g17641,
    g17642,g17644,g17645,I18609,g17648,I18614,g17651,g17652,g17672,g17673,I18647,g17676,
    g17677,I18653,g17680,g17681,g17683,g17684,I18662,g17687,I18667,I18674,g17691,g17707,
    g17709,g17710,I18694,g17713,g17714,I18700,g17717,g17718,g17720,g17721,I18709,g17733,
    g17735,g17737,g17738,I18728,g17741,g17742,I18734,g17745,g17746,g17754,g17756,g17758,
    g17759,I18752,g17762,g17763,I18758,g17772,g17774,g17776,g17777,I18778,I18788,g17782,
    I18795,g17789,g17791,g17794,g17811,I18810,g17812,I18813,g17815,I18822,g17818,I18825,
    I18829,g17821,I18832,g17844,I18835,I18839,g17847,I18842,g17870,I18845,I18849,g17873,
    I18852,g17926,I18855,g17929,I18858,g17952,I18861,g17953,I18865,g17955,I18868,g18008,
    g18061,I18872,g18062,I18875,g18065,g18088,I18879,g18091,I18882,I18885,g18093,I18888,
    I18891,I18894,I18897,I18900,I18903,I18906,I18909,I18912,g18102,I19012,g18200,I19235,
    g18421,I19238,g18422,I19345,g18527,I19348,g18528,I19384,g18562,I19484,g18660,I19487,
    g18661,g18827,g18828,g18829,g18830,g18831,g18832,I19661,g18833,g18874,g18875,g18876,
    g18877,g18878,g18880,I19671,I19674,g18882,g18883,g18884,g18885,g18886,g18887,g18888,
    g18889,g18891,g18892,g18894,g18895,g18896,g18897,g18898,g18903,g18904,g18905,g18907,
    g18908,g18911,g18916,g18917,I19704,g18918,I19707,g18926,g18929,g18930,g18931,g18932,
    g18938,g18939,I19719,g18940,g18944,g18945,g18946,g18947,g18948,g18952,g18953,g18954,
    I19734,g18957,g18975,g18976,g18977,g18978,g18979,g18980,g18983,g18984,g18988,g18989,
    g18990,g18991,I19756,g18997,I19759,g19050,I19762,g19061,g19067,g19068,g19071,I19772,
    g19074,I19775,g19127,I19778,g19128,g19144,g19146,I19786,g19147,I19789,g19200,g19208,
    I19796,g19210,I19799,g19263,I19802,g19264,g19273,g19276,I19813,g19277,g19330,I19818,
    g19343,g19345,g19351,g19352,I19831,g19353,g19355,I19837,g19360,I19843,g19361,g19362,
    g19364,g19365,g19366,I19851,g19367,g19368,g19369,g19370,I19857,g19371,g19373,g19374,
    I19863,g19375,g19376,g19379,g19385,g19386,g19387,g19389,g19394,g19395,g19396,g19397,
    g19398,g19399,g19407,g19408,g19409,g19410,g19411,g19412,g19414,g19415,g19416,g19417,
    g19421,g19427,g19428,g19429,g19431,g19432,g19433,g19434,g19435,g19437,g19438,g19439,
    g19440,g19443,g19445,I19917,g19446,g19451,g19452,g19454,I19927,g19458,g19468,g19469,
    g19470,g19471,g19472,g19473,g19476,g19477,g19478,g19479,g19480,g19481,g19482,g19489,
    g19490,g19491,g19492,g19493,g19494,g19498,g19499,g19502,g19503,g19504,g19505,g19517,
    g19518,g19519,g19520,g19523,g19524,g19526,g19527,g19528,g19529,g19531,g19532,g19533,
    g19537,g19538,g19539,g19541,g19542,g19543,g19544,g19552,g19553,g19554,g19558,g19559,
    g19565,g19566,g19567,g19569,g19570,g19573,g19574,g19577,g19579,g19580,g19586,I20035,
    g19592,g19600,g19602,g19603,g19606,g19609,g19612,g19617,g19618,g19620,g19626,g19629,
    g19630,g19633,g19634,g19635,g19636,g19638,g19644,g19649,g19650,g19652,g19653,g19654,
    g19657,g19658,g19659,g19662,g19666,g19670,g19672,g19673,g19675,g19676,g19677,g19678,
    g19679,g19682,g19683,g19685,g19686,g19687,g19688,g19689,g19690,g19694,g19695,g19696,
    g19697,g19698,I20116,g19699,g19709,g19710,g19711,g19712,g19713,g19714,g19718,g19719,
    I20130,g19720,g19730,g19731,g19732,g19733,g19734,g19737,g19738,g19739,g19741,g19742,
    g19743,g19744,g19745,g19747,g19748,g19750,g19751,g19753,g19754,g19755,g19757,g19760,
    g19761,g19762,g19763,g19765,g19766,g19769,g19770,g19771,g19772,g19773,g19776,g19777,
    g19779,g19780,g19781,g19783,g19785,g19786,g19787,g19789,g19790,g19794,g19798,g19799,
    g19800,I20216,g19801,g19852,g19860,g19861,I20233,g19862,g19865,g19866,g19869,g19872,
    g19878,g19881,g19882,g19885,g19902,g19905,g19908,g19912,g19915,g19930,g19931,g19947,
    g19950,g19952,g19954,g19957,g19960,g19961,g19963,g19964,g19979,g19980,g19996,g19998,
    g20004,g20005,g20006,g20008,g20009,g20010,g20025,g20026,g20028,g20033,g20035,g20036,
    g20037,g20038,g20040,g20041,g20046,I20318,I20321,g20050,g20052,g20053,g20054,g20057,
    g20058,g20059,g20060,g20064,g20065,g20066,g20067,g20070,g20071,g20072,g20073,g20078,
    g20079,g20080,g20085,I20355,g20086,g20087,g20088,g20089,g20090,g20091,g20096,g20097,
    I20369,g20100,g20101,g20102,g20103,g20104,g20105,g20106,g20110,g20113,I20385,g20114,
    I20388,g20127,g20128,g20129,g20130,g20132,I20399,g20136,g20144,g20145,g20146,g20147,
    g20153,I20412,g20154,g20157,g20158,g20159,g20164,g20166,g20167,g20168,I20433,g20175,
    g20178,g20179,g20180,g20182,I20447,g20189,g20190,g20191,g20192,g20194,g20195,g20197,
    g20204,g20207,g20208,g20209,g20210,g20211,g20212,g20213,I20495,g20219,g20229,I20499,
    g20230,g20231,g20232,g20233,g20235,g20237,g20238,g20239,g20240,g20242,g20247,g20265,
    g20266,g20267,g20268,g20269,g20270,g20272,g20273,g20274,g20275,g20277,I20529,g20283,
    g20320,g20321,g20322,g20323,g20324,g20325,g20326,g20327,g20328,g20329,I20542,g20330,
    g20372,g20373,g20374,g20379,g20380,g20381,g20382,g20383,g20384,g20385,g20386,g20387,
    g20388,g20389,I20562,g20391,g20432,g20433,g20434,g20435,I20569,g20436,g20441,g20442,
    g20443,g20444,g20445,g20446,g20447,g20448,g20449,g20450,g20451,g20452,I20584,g20453,
    g20494,g20495,g20496,g20497,g20498,g20499,g20500,g20501,g20502,g20503,g20504,g20505,
    g20506,g20507,g20508,g20509,g20510,g20511,g20512,g20513,g20514,g20515,I20609,g20516,
    g20523,g20524,g20525,g20526,g20527,g20528,g20529,g20530,g20531,g20532,g20533,g20534,
    g20535,g20536,g20537,g20538,g20539,g20540,g20541,g20542,g20543,g20544,g20545,g20546,
    g20547,g20548,g20549,g20550,g20551,g20552,g20553,g20554,g20555,g20556,I20647,I20650,
    g20558,g20560,g20561,g20562,g20563,g20564,g20565,g20566,g20567,g20568,g20569,g20570,
    g20571,g20572,g20573,g20574,g20575,g20576,g20577,g20578,g20579,g20580,g20582,g20583,
    g20584,g20585,g20586,g20587,g20588,g20589,g20590,g20591,g20592,g20593,g20594,g20595,
    I20690,g20596,g20597,g20598,g20599,g20600,g20601,g20603,g20604,g20605,g20606,g20607,
    g20608,g20609,g20610,g20611,g20612,g20613,g20614,g20615,g20616,g20617,g20618,g20622,
    g20623,g20624,g20625,g20626,g20627,g20629,g20630,g20631,g20632,g20633,g20634,g20635,
    g20636,g20637,g20638,g20639,g20640,g20641,g20642,g20643,g20648,g20649,g20650,g20651,
    I20744,I20747,g20653,I20750,I20753,g20655,g20656,g20657,g20659,g20660,g20661,g20662,
    g20663,g20664,g20665,g20666,g20667,g20668,g20669,g20670,g20671,g20672,g20673,g20674,
    g20679,g20680,g20681,I20781,g20695,g20696,g20697,g20698,g20699,g20700,g20701,g20702,
    g20703,g20704,I20793,g20705,g20706,g20707,g20708,g20709,g20710,g20711,g20712,g20713,
    g20714,g20715,g20716,g20732,g20737,g20738,I20816,I20819,g20764,g20765,g20766,g20767,
    g20768,g20769,g20770,g20771,g20772,I20830,g20773,g20774,g20775,g20776,g20777,g20778,
    g20779,g20780,I20840,g20781,g20782,I20846,g20785,g20852,g20853,g20869,g20874,I20861,
    I20864,g20900,I20867,I20870,g20902,g20903,g20904,g20909,g20910,g20911,g20912,g20913,
    g20914,I20882,g20915,g20916,g20917,g20918,g20919,g20920,g20921,I20891,g20922,g20923,
    I20895,g20924,g20978,g20993,g20994,g21010,I20910,g21036,I20913,g21037,g21048,g21049,
    g21050,g21051,g21052,g21053,g21054,g21055,g21056,g21057,g21058,g21059,g21060,I20929,
    g21061,g21068,g21069,I20937,g21070,g21123,g21138,g21139,g21155,g21156,g21160,I20951,
    g21175,I20954,I20957,g21177,g21178,g21179,g21180,g21181,g21182,g21183,g21184,g21185,
    g21189,g21204,g21205,g21221,g21222,g21225,g21228,I20982,I20985,g21246,g21247,g21248,
    g21249,g21252,g21267,g21268,g21269,I20999,I21002,g21271,I21006,g21273,g21274,g21275,
    I21013,g21278,g21279,g21280,g21281,I21019,g21282,g21286,I21029,g21290,g21291,I21033,
    I21036,g21293,g21295,I21042,g21297,g21299,I21047,g21300,g21304,g21305,g21306,g21308,
    I21058,g21326,g21329,I21067,g21335,g21336,g21337,I21074,g21340,g21343,g21346,g21349,
    g21352,g21355,g21358,g21362,I21100,g21366,g21369,g21370,g21379,g21380,g21381,g21383,
    I21115,g21387,g21393,g21395,g21396,g21397,g21398,g21399,g21400,g21406,g21407,g21408,
    g21409,g21410,g21411,g21412,g21413,g21414,g21418,g21421,g21422,g21423,g21424,g21425,
    g21426,g21427,g21428,g21430,g21431,g21434,I21162,g21451,g21454,g21455,g21456,g21457,
    g21458,g21460,g21461,g21463,g21466,g21467,I21181,g21468,g21510,g21511,I21189,g21514,
    g21556,g21560,g21561,I21199,g21562,g21604,g21607,g21608,g21609,g21610,I21210,g21611,
    g21653,g21654,g21656,g21657,g21659,g21660,I21222,g21661,g21662,I21226,g21665,g21666,
    I21230,g21669,g21670,I21234,g21673,g21674,I21238,g21677,g21678,I21242,g21681,g21682,
    I21246,g21685,g21686,I21250,g21689,g21690,I21254,g21693,g21694,I21258,g21697,I21285,
    g21722,I21288,g21723,I21291,g21724,I21294,g21725,I21297,g21726,I21300,I21477,g21902,
    I21480,g21903,I21483,g21904,I21486,g21905,g22136,g22137,g22138,I21722,g22139,g22144,
    g22146,g22147,g22148,g22150,I21734,g22151,g22153,g22154,g22155,g22156,I21744,g22159,
    g22166,g22167,g22168,g22169,g22170,g22171,I21757,g22173,g22176,g22177,g22178,g22179,
    g22180,g22181,I21766,g22182,I21769,g22189,g22192,I21776,g22194,g22197,g22198,g22199,
    g22200,g22201,I21784,g22202,I21787,g22207,I21792,g22210,g22213,g22214,g22215,I21802,
    g22220,g22223,g22224,g22227,I21810,g22228,I21815,g22300,g22303,g22305,g22311,g22317,
    I21831,g22319,g22330,I21838,g22332,g22338,g22339,g22341,g22358,g22359,I21849,g22360,
    g22406,g22407,g22408,I21860,g22409,g22449,g22455,g22456,g22492,g22493,g22494,g22495,
    g22496,g22497,g22519,g22520,g22526,g22527,g22528,g22529,I21911,g22541,g22542,g22543,
    g22544,I21918,g22546,I21922,g22550,I21930,g22592,g22593,I21934,g22594,I21941,g22626,
    g22635,g22646,I21959,g22647,g22649,I21969,g22658,g22660,g22667,g22682,I22000,g22683,
    I22009,g22698,g22714,g22716,g22718,I22024,g22719,I22028,g22721,I22031,g22722,g22756,
    g22758,g22759,g22761,I22046,g22763,g22830,g22840,g22841,g22842,g22844,g22845,g22847,
    g22854,g22855,g22856,g22857,g22858,g22860,g22865,g22866,g22867,g22868,g22869,g22870,
    I22096,g22881,g22882,g22883,g22884,g22896,g22897,g22898,g22903,I22111,g22904,I22114,
    g22905,g22906,g22907,g22919,g22922,I22124,g22923,g22926,I22128,g22927,I22131,g22928,
    g22935,g22936,I22143,g22957,g22973,g22974,g22975,I22149,g22976,g22979,I22153,g22980,
    g22981,g22985,g22986,g22987,g22988,g22989,g22994,g22995,g22996,g22997,g22998,g22999,
    g23000,g23001,I22177,I22180,g23003,g23004,g23005,g23011,g23012,g23013,g23014,g23015,
    g23016,g23017,g23018,g23019,g23020,g23021,g23022,g23026,g23027,g23028,g23029,g23030,
    g23031,I22211,g23032,g23041,g23046,g23055,g23057,g23058,g23059,g23060,g23061,g23066,
    g23082,g23084,g23085,g23086,I22240,g23088,g23111,g23127,g23128,g23138,g23152,I22264,
    g23154,g23170,I22275,g23172,g23182,g23189,I22286,I22289,g23191,g23192,g23196,I22302,
    g23202,g23203,g23211,g23214,g23215,g23216,I22316,g23219,g23221,g23222,g23223,g23226,
    g23227,g23228,I22327,g23230,g23231,I22331,g23232,g23233,g23234,g23235,g23236,g23237,
    g23238,g23239,g23242,g23243,I22343,g23244,g23245,g23246,g23247,g23248,g23249,g23250,
    I22353,g23252,g23253,g23256,g23257,g23258,g23259,g23260,I22366,g23263,g23264,g23267,
    g23270,g23271,g23272,g23273,g23274,I22380,g23277,g23278,g23279,g23282,g23283,g23284,
    g23285,g23289,g23290,g23291,I22400,g23299,g23300,g23301,g23302,g23303,g23304,g23305,
    g23306,g23307,g23308,g23312,g23313,I22419,g23320,I22422,g23321,I22425,g23322,g23323,
    g23331,g23332,g23333,g23334,g23335,g23336,g23337,g23338,g23339,g23340,g23341,I22444,
    g23347,g23350,g23351,g23352,g23353,g23354,g23355,g23356,I22458,g23359,I22461,g23360,
    I22464,g23361,I22467,g23362,I22470,g23363,g23375,g23376,g23377,g23378,g23380,g23382,
    I22485,g23384,I22488,g23385,g23388,g23390,g23391,g23393,I22499,g23394,I22502,g23395,
    g23398,g23399,g23400,g23402,I22512,g23403,g23406,g23408,g23409,g23410,g23411,g23413,
    I22525,g23414,g23417,g23418,g23419,g23420,g23421,g23422,g23423,g23425,I22539,g23426,
    I22542,g23427,g23429,I22547,g23430,g23431,g23432,g23433,g23434,g23435,I22557,g23440,
    g23443,I22561,g23444,I22564,g23445,g23446,g23447,g23448,g23449,I22571,g23450,g23452,
    I22576,g23453,g23456,I22580,g23457,I22583,g23458,g23459,g23460,g23461,I22589,g23462,
    g23472,g23473,g23476,g23477,g23478,g23479,I22601,g23480,I22604,g23481,g23482,g23483,
    g23485,g23486,g23487,g23488,g23489,g23490,g23491,g23492,g23493,I22619,g23494,I22622,
    g23495,g23496,g23499,g23500,g23501,g23502,g23503,g23504,g23505,g23506,g23507,g23508,
    g23509,g23510,I22640,g23511,g23512,g23515,g23516,g23517,g23518,g23519,g23520,g23521,
    g23522,g23523,g23524,g23525,g23526,g23527,g23528,g23529,g23530,I22665,g23534,g23537,
    g23538,g23539,g23541,g23542,g23543,g23544,g23545,g23546,g23547,g23548,g23549,g23550,
    I22692,g23555,g23558,g23559,g23563,g23565,g23566,g23567,g23568,g23569,g23570,g23571,
    g23573,I22725,g23578,I22729,g23582,g23585,g23589,g23605,g23607,g23608,g23609,g23610,
    g23611,I22745,I22748,g23613,g23614,I22769,g23620,g23629,g23645,g23647,g23648,g23649,
    g23650,g23651,I22785,I22788,g23653,g23654,g23665,g23681,I22816,I22819,g23684,g23698,
    g23714,g23715,g23732,g23745,g23746,g23749,I22886,I22889,g23760,g23764,g23767,g23768,
    g23769,g23776,I22918,g23777,g23787,g23788,g23789,g23792,g23793,g23794,g23800,g23812,
    g23813,g23814,g23815,g23816,g23819,g23820,g23821,I22989,g23823,g23824,g23838,g23839,
    g23840,g23841,g23842,g23843,g23844,g23847,g23848,g23849,g23858,g23859,g23860,g23861,
    g23862,g23863,g23864,g23865,g23868,g23869,g23870,g23874,g23875,g23876,g23877,g23878,
    g23879,g23880,g23881,g23882,g23886,g23887,g23888,g23889,g23893,g23894,g23895,g23896,
    g23897,g23898,g23899,g23902,g23903,g23904,g23905,g23906,g23907,g23908,g23912,g23913,
    g23914,g23915,g23916,g23922,g23923,g23924,g23925,g23926,g23927,g23928,g23929,g23930,
    g23931,g23935,g23936,g23937,g23938,g23939,g23940,g23941,g23942,g23943,g23944,g23945,
    g23946,g23947,g23948,g23952,g23953,I23099,g23954,g23961,g23962,g23963,g23964,g23965,
    g23966,g23967,g23968,g23969,g23970,g23971,g23982,g23983,g23984,g23985,g23986,g23987,
    g23988,g23992,g23993,g23994,g23995,g23999,g24000,g24003,I23149,g24005,g24010,g24013,
    g24017,g24019,g24020,g24021,g24022,g24023,g24024,g24025,g24026,g24027,g24028,g24029,
    g24030,g24031,g24032,g24033,g24034,g24035,g24036,g24037,g24038,g24039,g24040,g24041,
    g24042,g24043,g24044,g24045,g24046,g24047,g24048,g24049,g24050,g24051,g24052,g24053,
    g24054,g24055,g24056,g24057,g24058,g24059,g24060,g24061,g24062,g24063,g24064,g24065,
    g24066,g24067,g24068,g24069,g24070,g24071,g24072,g24073,g24074,g24075,g24076,g24077,
    g24078,g24079,g24080,g24081,g24082,g24083,g24084,g24085,g24086,g24087,g24088,g24089,
    g24090,g24091,g24092,g24093,g24094,g24095,g24096,g24097,g24098,g24099,g24100,g24101,
    g24102,g24103,g24104,g24105,g24106,g24107,g24108,g24109,g24110,g24111,g24112,g24113,
    g24114,g24115,g24116,g24117,g24118,g24119,g24120,g24121,g24122,g24123,g24124,g24125,
    g24126,g24127,g24128,g24129,g24130,g24131,g24132,g24133,g24134,g24135,g24136,g24137,
    g24138,g24146,g24147,g24149,g24150,I23300,g24152,I23303,g24153,I23306,g24154,I23309,
    g24155,I23312,g24156,I23315,g24157,I23318,g24158,I23321,g24159,I23324,g24160,I23327,
    g24161,I23330,g24162,I23333,g24163,I23336,g24164,I23339,g24165,I23342,g24166,I23345,
    g24167,I23348,g24168,I23351,g24169,I23354,g24170,I23357,g24171,I23360,g24172,I23363,
    g24173,I23366,g24174,I23369,g24175,I23372,g24176,I23375,g24177,I23378,g24178,I23381,
    g24179,I23384,g24180,I23387,g24181,I23390,g24182,I23393,g24183,I23396,g24184,I23399,
    g24185,g24356,g24357,g24358,g24359,g24360,g24361,g24364,g24365,g24366,g24367,g24368,
    g24372,g24373,g24375,g24376,g24377,g24379,g24384,g24385,g24386,g24388,g24389,g24394,
    g24396,g24397,g24404,g24405,g24407,g24417,g24418,g24419,g24424,g24425,g24426,g24428,
    g24429,g24431,g24437,g24438,g24452,g24463,I23671,g24466,g24474,I23680,g24477,I23684,
    g24481,I23688,g24483,I23694,g24489,g24490,g24505,I23711,g24506,g24509,g24515,g24516,
    g24522,g24524,g24525,g24526,g24527,g24533,g24534,g24535,g24540,g24548,g24560,g24568,
    g24571,g24579,g24585,g24586,g24587,g24603,g24604,g24605,g24623,g24625,g24626,g24636,
    g24648,g24655,g24665,g24667,g24683,g24685,g24699,g24711,g24718,g24732,g24744,g24756,
    g24759,g24770,g24778,g24789,g24791,g24795,g24818,I23998,g24819,g24825,I24008,g24836,
    g24839,I24022,g24850,I24038,g24866,I24041,g24869,g24891,I24060,g24893,I24078,g24911,
    I24089,g24920,g24960,g24963,I24128,g24964,g24966,g24971,g24978,g24979,g24980,g24981,
    g24982,g24985,g24986,g24987,g24991,g24992,g24993,g24994,g24995,g24996,g24999,g25000,
    g25001,g25006,g25007,g25008,g25009,g25011,g25013,g25015,g25016,g25017,g25023,g25024,
    g25025,I24191,g25027,g25032,g25034,g25035,g25036,g25039,g25044,g25046,g25047,I24215,
    g25051,g25055,g25060,I24228,g25064,g25070,g25072,I24237,g25073,g25080,g25081,g25082,
    g25083,g25090,g25092,g25097,g25098,g25099,g25100,g25101,g25109,g25111,I24278,I24281,
    g25115,g25116,g25117,g25118,g25119,g25120,g25121,g25131,g25133,g25134,g25135,g25136,
    g25137,g25138,g25139,g25140,g25153,g25154,g25155,g25156,g25157,g25158,I24331,I24334,
    g25168,g25169,g25170,g25171,g25174,g25180,g25182,g25183,g25184,g25185,g25188,g25193,
    g25194,g25195,g25196,g25197,g25198,g25202,g25206,g25208,g25209,g25210,g25211,g25212,
    g25213,g25214,g25218,I24393,I24396,g25220,g25221,I24400,g25222,g25224,g25225,g25226,
    g25227,g25228,g25230,g25231,g25232,g25239,g25240,g25241,g25242,g25243,g25244,g25245,
    g25246,g25248,g25249,I24434,g25250,I24445,I24448,g25260,g25262,g25263,g25264,I24455,
    g25265,g25266,g25267,g25272,g25273,g25274,g25282,g25283,I24474,g25284,g25286,g25287,
    g25288,g25289,g25296,g25297,g25298,g25299,g25307,g25308,g25316,I24497,g25322,g25324,
    g25325,g25326,g25327,g25340,g25348,g25356,g25369,g25370,g25380,g25388,g25399,g25409,
    g25410,I24558,g25423,g25424,g25438,g25451,g25452,g25465,g25480,g25481,g25505,g25506,
    g25513,g25517,g25523,g25524,g25525,g25528,g25529,g25533,g25534,g25535,g25538,g25541,
    g25542,g25544,g25546,g25547,g25548,g25549,g25550,g25552,g25553,g25554,g25555,g25556,
    g25557,g25558,g25560,g25561,g25562,g25563,g25564,g25566,I24759,g25620,I24781,g25640,
    I24784,g25641,I24787,g25642,I24839,g25692,g25766,I24920,g25771,g25773,g25781,g25783,
    g25786,g25790,g25820,g25830,g25837,g25838,g25849,g25869,g25882,g25886,g25892,g25893,
    g25899,I25005,g25903,I25028,g25930,g25994,I25095,g25997,I25105,g26026,g26054,I25115,
    g26055,g26081,g26083,g26093,I25146,g26105,I25161,g26131,I25190,g26187,g26260,g26284,
    g26326,g26337,g26340,I25327,g26364,I25351,g26400,I25356,g26424,I25359,g26483,I25366,
    g26488,I25369,g26510,g26518,I25380,g26519,g26548,I25391,g26549,g26575,I25399,g26576,
    g26605,g26607,g26608,g26614,g26615,g26631,g26632,g26634,g26648,g26653,g26654,g26655,
    g26656,g26672,g26679,g26680,g26681,g26682,g26683,g26693,g26700,g26701,g26702,g26709,
    g26710,g26718,g26720,g26724,g26731,g26732,g26736,g26743,g26744,g26754,g26758,g26765,
    g26769,g26776,g26777,g26784,g26788,g26792,I25511,I25514,g26802,g26803,g26804,g26810,
    g26811,g26812,g26814,g26816,g26817,I25530,g26818,I25534,g26820,g26824,I25541,g26825,
    g26827,g26830,g26831,g26832,I25552,g26834,I25555,g26835,g26836,g26837,I25562,g26840,
    g26841,I25567,g26843,I25576,g26850,I25579,g26851,I25586,g26856,I25591,g26859,I25594,
    g26860,I25598,g26862,g26869,I25606,g26870,I25677,g26935,I25680,g26936,I25683,g26937,
    I25689,g26941,I25692,g26942,I25695,g26943,g26973,g26987,g26990,g27004,g27009,g27011,
    I25743,g27013,g27014,g27015,g27017,I25750,g27018,g27038,I25779,g27051,I25786,g27064,
    I25790,g27074,g27084,g27088,g27089,g27091,g27092,g27100,g27101,g27112,g27142,g27155,
    I25869,g27163,I25882,g27187,g27237,g27242,g27245,g27279,I26004,g27320,g27349,I26100,
    g27402,g27415,I26130,g27438,g27492,I26195,g27527,g27554,g27565,g27573,g27576,g27583,
    g27585,g27592,g27597,I26296,g27662,I26309,g27675,g27698,I26334,g27708,I26337,g27709,
    g27730,I26356,g27736,g27737,I26378,g27773,I26381,g27774,g27830,I26406,I26409,g27832,
    I26427,g27880,I26430,g27881,g27928,I26448,g27929,I26451,g27930,I26466,g27956,g27961,
    I26479,g27967,g27971,g27975,g27976,g27977,g27983,g27984,g27985,g27989,g27990,g27991,
    I26503,g27993,g27994,I26508,g27996,I26512,g27998,I26516,g28009,g28032,g28033,g28034,
    g28036,g28037,g28038,g28039,g28040,I26578,g28079,I26581,g28080,I26584,g28081,g28119,
    g28120,g28121,g28126,g28127,I26638,g28137,I26649,g28142,I26654,g28147,I26664,g28155,
    I26667,g28156,I26670,g28157,I26676,g28161,I26679,g28162,I26682,g28163,I26687,g28166,
    I26693,g28173,I26700,g28181,I26705,g28184,I26710,g28187,g28241,g28250,I26785,g28262,
    I26799,g28274,g28294,g28307,g28321,g28325,g28326,I26880,g28367,g28370,g28380,g28399,
    I26925,g28431,I26929,g28436,g28441,I26936,g28443,I26952,g28463,g28479,I26989,g28508,
    g28559,g28575,g28579,g28590,g28593,g28598,g28604,g28606,g28608,g28615,g28620,g28633,
    g28648,g28656,g28669,g28675,g28678,g28693,g28696,I27192,g28709,g28711,g28713,g28726,
    I27232,g28752,I27235,I27238,g28754,I27253,g28779,I27271,g28819,I27314,g28917,g28918,
    g28954,I27368,g29013,g29014,I27385,g29041,I27388,g29042,I27391,g29043,g29044,g29045,
    g29056,I27401,g29067,g29079,g29080,g29081,g29092,g29093,g29115,g29116,g29117,g29128,
    g29129,g29130,I27449,g29147,g29149,g29150,g29151,g29152,g29153,g29169,g29170,g29171,
    g29172,g29177,I27481,g29185,g29190,I27492,g29194,I27495,g29195,g29196,I27543,g29209,
    I27546,I27549,I27552,I27555,I27558,I27561,I27564,I27567,I27570,I27573,I27576,I27579,
    g29310,g29311,g29312,I27677,g29317,g29318,g29333,g29339,g29342,g29343,g29348,I27713,
    g29353,I27718,g29358,g29365,I27730,g29368,I27735,g29371,I27738,g29372,I27742,g29374,
    I27749,g29379,g29385,I27758,g29474,I27777,g29491,I27784,g29498,g29505,g29507,g29597,
    I27927,g29653,I27941,g29669,I27954,g29689,g29697,g29707,I27970,g29713,g29725,g29744,
    g29745,I28002,g29755,I28014,g29765,g29800,g29811,g29812,I28062,g29814,g29846,g29847,
    g29862,g29863,g29878,g29893,I28128,g29897,g29905,g29906,g29911,g29912,g29913,g29920,
    g29921,g29922,g29923,g29925,g29927,g29928,g29929,I28162,g29930,g29939,g29941,g29942,
    g29944,I28174,g29945,g29948,g29950,g29953,g29955,I28185,g29956,g29960,g29961,g29963,
    g29965,g29967,I28199,g29970,g29976,g29977,g29978,g29980,g29981,g29983,g29993,g29994,
    g29995,g29996,g29997,g29998,g29999,I28241,g30012,g30016,g30017,g30018,g30019,g30020,
    g30021,g30022,g30036,g30037,g30038,g30039,g30040,g30052,g30053,g30054,g30055,g30063,
    g30065,g30067,g30068,I28301,g30072,g30074,g30076,g30077,g30079,g30085,g30087,g30088,
    g30090,g30097,g30100,g30102,I28336,g30105,g30113,I28349,g30116,g30142,I28390,g30155,
    I28419,g30182,g30184,I28434,g30195,g30206,I28458,g30217,g30218,I28480,g30237,g30259,
    g30292,I28540,g30295,g30296,g30297,g30299,I28548,g30301,g30302,g30303,g30305,g30306,
    g30309,g30310,g30312,g30313,g30318,I28572,g30321,g30322,I28576,g30325,I28579,g30326,
    I28582,I28585,g30328,I28588,I28591,I28594,I28597,I28832,g30565,g30567,g30568,I28838,
    g30569,g30572,g30578,I28851,g30591,g30593,I28866,g30606,I28872,g30610,I28883,g30729,
    I28897,g30917,I28908,g30928,I28913,g30931,g30983,g30989,g30990,I28925,g30991,g30996,
    g30997,g30998,g30999,g31000,g31013,g31138,I29002,g31189,I29013,g31213,g31227,g31239,
    g31243,I29139,g31479,I29149,g31487,I29182,I29185,g31522,I29199,g31578,I29204,g31596,
    I29207,g31601,g31608,I29211,g31609,I29214,g31616,g31623,I29218,g31624,I29221,g31631,
    g31638,I29225,g31639,I29228,g31646,g31653,I29233,g31655,I29236,I29239,g31657,I29242,
    g31658,I29245,I29248,g31666,g31667,I29337,g31771,I29363,g31791,I29368,g31794,I29371,
    g31795,g31796,g31797,g31798,g31799,g31800,g31801,g31802,g31803,g31804,g31805,g31806,
    g31807,g31808,g31809,g31810,g31811,g31812,g31813,g31814,g31815,g31816,g31817,g31818,
    g31819,g31820,g31821,g31822,g31823,g31824,g31825,g31826,g31827,g31828,g31829,g31830,
    g31831,g31832,g31833,g31834,g31835,g31836,g31837,g31838,g31839,g31840,g31841,g31842,
    g31843,g31844,g31845,g31846,g31847,g31848,g31849,g31850,g31851,g31852,g31853,g31854,
    g31855,g31856,g31857,g31858,g31859,I29438,I29441,I29444,I29447,g31937,g31945,I29571,
    g32015,I29579,g32021,I29582,g32024,I29585,g32027,g32033,g32038,g32090,g32099,g32118,
    g32137,g32138,I29717,I29720,g32186,g32192,g32201,g32318,g32329,I29891,g32363,I29894,
    g32364,g32377,I29909,g32381,g32382,I29913,g32383,g32384,g32393,g32394,I29936,g32404,
    I29939,g32407,g32415,g32421,g32430,I29961,g32433,g32434,I29965,g32437,g32438,I29969,
    g32441,g32442,I29973,g32445,g32446,I29977,g32449,g32450,I29981,g32453,g32456,g32457,
    g32458,g32459,g32460,g32461,g32462,g32463,g32464,g32465,g32466,g32467,g32468,g32469,
    g32470,g32471,g32472,g32473,g32474,g32475,g32476,g32477,g32478,g32479,g32480,g32481,
    g32482,g32483,g32484,g32485,g32486,g32487,g32488,g32489,g32490,g32491,g32492,g32493,
    g32494,g32495,g32496,g32497,g32498,g32499,g32500,g32501,g32502,g32503,g32504,g32505,
    g32506,g32507,g32508,g32509,g32510,g32511,g32512,g32513,g32514,g32515,g32516,g32517,
    g32518,g32519,g32521,g32522,g32523,g32524,g32525,g32526,g32527,g32528,g32529,g32530,
    g32531,g32532,g32533,g32534,g32535,g32536,g32537,g32538,g32539,g32540,g32541,g32542,
    g32543,g32544,g32545,g32546,g32547,g32548,g32549,g32550,g32551,g32552,g32553,g32554,
    g32555,g32556,g32557,g32558,g32559,g32560,g32561,g32562,g32563,g32564,g32565,g32566,
    g32567,g32568,g32569,g32570,g32571,g32572,g32573,g32574,g32575,g32576,g32577,g32578,
    g32579,g32580,g32581,g32582,g32583,g32584,g32586,g32587,g32588,g32589,g32590,g32591,
    g32592,g32593,g32594,g32595,g32596,g32597,g32598,g32599,g32600,g32601,g32602,g32603,
    g32604,g32605,g32606,g32607,g32608,g32609,g32610,g32611,g32612,g32613,g32614,g32615,
    g32616,g32617,g32618,g32619,g32620,g32621,g32622,g32623,g32624,g32625,g32626,g32627,
    g32628,g32629,g32630,g32631,g32632,g32633,g32634,g32635,g32636,g32637,g32638,g32639,
    g32640,g32641,g32642,g32643,g32644,g32645,g32646,g32647,g32648,g32649,g32651,g32652,
    g32653,g32654,g32655,g32656,g32657,g32658,g32659,g32660,g32661,g32662,g32663,g32664,
    g32665,g32666,g32667,g32668,g32669,g32670,g32671,g32672,g32673,g32674,g32675,g32676,
    g32677,g32678,g32679,g32680,g32681,g32682,g32683,g32684,g32685,g32686,g32687,g32688,
    g32689,g32690,g32691,g32692,g32693,g32694,g32695,g32696,g32697,g32698,g32699,g32700,
    g32701,g32702,g32703,g32704,g32705,g32706,g32707,g32708,g32709,g32710,g32711,g32712,
    g32713,g32714,g32716,g32717,g32718,g32719,g32720,g32721,g32722,g32723,g32724,g32725,
    g32726,g32727,g32728,g32729,g32730,g32731,g32732,g32733,g32734,g32735,g32736,g32737,
    g32738,g32739,g32740,g32741,g32742,g32743,g32744,g32745,g32746,g32747,g32748,g32749,
    g32750,g32751,g32752,g32753,g32754,g32755,g32756,g32757,g32758,g32759,g32760,g32761,
    g32762,g32763,g32764,g32765,g32766,g32767,g32768,g32769,g32770,g32771,g32772,g32773,
    g32774,g32775,g32776,g32777,g32778,g32779,g32781,g32782,g32783,g32784,g32785,g32786,
    g32787,g32788,g32789,g32790,g32791,g32792,g32793,g32794,g32795,g32796,g32797,g32798,
    g32799,g32800,g32801,g32802,g32803,g32804,g32805,g32806,g32807,g32808,g32809,g32810,
    g32811,g32812,g32813,g32814,g32815,g32816,g32817,g32818,g32819,g32820,g32821,g32822,
    g32823,g32824,g32825,g32826,g32827,g32828,g32829,g32830,g32831,g32832,g32833,g32834,
    g32835,g32836,g32837,g32838,g32839,g32840,g32841,g32842,g32843,g32844,g32846,g32847,
    g32848,g32849,g32850,g32851,g32852,g32853,g32854,g32855,g32856,g32857,g32858,g32859,
    g32860,g32861,g32862,g32863,g32864,g32865,g32866,g32867,g32868,g32869,g32870,g32871,
    g32872,g32873,g32874,g32875,g32876,g32877,g32878,g32879,g32880,g32881,g32882,g32883,
    g32884,g32885,g32886,g32887,g32888,g32889,g32890,g32891,g32892,g32893,g32894,g32895,
    g32896,g32897,g32898,g32899,g32900,g32901,g32902,g32903,g32904,g32905,g32906,g32907,
    g32908,g32909,g32911,g32912,g32913,g32914,g32915,g32916,g32917,g32918,g32919,g32920,
    g32921,g32922,g32923,g32924,g32925,g32926,g32927,g32928,g32929,g32930,g32931,g32932,
    g32933,g32934,g32935,g32936,g32937,g32938,g32939,g32940,g32941,g32942,g32943,g32944,
    g32945,g32946,g32947,g32948,g32949,g32950,g32951,g32952,g32953,g32954,g32955,g32956,
    g32957,g32958,g32959,g32960,g32961,g32962,g32963,g32964,g32965,g32966,g32967,g32968,
    g32969,g32970,g32971,g32972,g32973,g32974,I30537,g33072,I30641,I30644,g33080,I30686,
    g33120,g33127,g33136,g33142,I30766,g33228,g33246,g33250,g33258,g33326,I30861,g33335,
    g33346,g33354,g33375,I30901,g33377,I30904,g33378,g33382,g33385,g33388,g33391,g33413,
    g33424,g33426,g33430,I30959,I30962,g33436,g33442,I30971,g33443,g33451,I30980,g33454,
    I30983,g33455,I30986,g33456,I30989,g33457,I30992,g33458,I30995,g33459,I30998,g33460,
    I31361,I31459,g33631,g33635,I31463,I31466,g33637,I31469,g33638,I31474,g33641,I31477,
    g33645,I31482,g33648,I31486,g33653,g33658,I31491,I31494,g33660,I31497,g33661,I31500,
    g33665,I31504,g33670,I31515,g33682,g33686,I31523,g33688,I31528,g33691,g33695,I31535,
    g33696,I31539,g33698,I31545,g33702,I31550,g33705,I31555,g33708,I31561,g33712,I31564,
    g33713,I31569,g33716,I31581,g33726,I31586,g33729,I31597,g33736,I31604,g33744,I31607,
    g33750,I31610,g33755,I31616,g33761,I31619,g33766,I31622,g33772,I31625,g33778,g33797,
    g33799,I31642,g33800,g33804,I31650,g33806,I31659,g33813,I31672,g33827,I31686,g33839,
    I31694,g33845,I31701,g33850,I31724,I31727,g33875,g33888,I31748,I31751,g33895,I31770,
    g33912,I31776,g33916,I31779,g33917,I31782,g33918,I31786,g33920,I31791,g33923,I31796,
    g33926,I31800,g33928,I31803,g33929,I31807,g33931,I31810,g33932,I31814,g33934,I31817,
    I31820,g33936,I31823,g33937,I31829,g33944,I31878,g34042,g34044,g34047,g34049,g34052,
    g34053,g34058,g34059,g34060,g34062,g34068,g34070,g34094,I32051,g34118,I32056,g34121,
    I32059,g34122,I32062,g34123,g34124,I32067,g34126,I32071,g34130,I32074,g34131,g34132,
    I32079,g34134,I32089,g34142,I32093,g34144,I32096,g34145,g34147,I32103,g34150,I32106,
    g34151,I32109,g34152,g34156,I32116,g34159,I32119,g34160,g34161,g34181,g34188,g34192,
    I32150,g34195,g34197,g34200,I32158,I32161,g34202,g34208,I32170,g34209,I32173,g34210,
    I32192,I32195,g34222,g34229,I32222,g34241,I32225,g34242,I32228,g34243,I32231,g34244,
    I32234,g34245,I32237,g34246,I32240,g34247,I32243,g34248,g34270,g34271,g34272,g34275,
    g34276,I32274,g34277,I32284,g34285,I32297,g34296,g34299,I32305,g34302,I32309,g34304,
    g34307,g34308,g34311,g34312,g34313,g34315,g34316,g34317,g34320,g34323,g34325,g34326,
    g34327,g34328,g34336,g34339,g34343,I32352,g34345,g34346,g34351,I32364,g34358,I32388,
    I32391,g34384,g34387,g34391,g34392,g34400,g34408,g34409,g34418,g34419,g34420,g34423,
    I32446,I32449,g34426,I32452,g34427,I32455,g34428,I32458,g34429,I32461,g34430,I32464,
    g34431,I32467,g34432,I32470,g34433,I32473,g34434,I32476,I32479,I32482,g34471,I32525,
    g34472,g34473,I32535,g34480,I32547,g34490,I32550,g34491,g34501,g34504,g34505,g34510,
    g34511,g34512,g34521,g34522,I32591,g34530,I32594,g34531,I32601,g34536,g34539,I32607,
    g34540,g34543,I32613,g34544,I32617,g34549,I32621,g34553,g34559,I32639,g34569,g34570,
    I32645,g34573,I32648,g34574,I32651,g34575,I32654,g34576,I32659,g34579,I32665,g34583,
    I32671,g34587,I32675,g34589,I32678,g34590,I32681,g34591,I32684,g34592,I32687,g34593,
    I32690,g34594,I32693,g34595,I32696,g34596,I32699,I32752,g34648,I32763,g34653,I32766,
    g34654,I32770,g34656,I32775,g34659,g34660,I32782,g34664,I32788,g34668,I32791,g34669,
    I32794,g34670,I32797,g34671,I32800,g34672,I32803,g34673,I32806,g34674,I32809,g34675,
    I32812,g34676,I32815,g34677,I32820,g34680,I32824,g34682,I32827,g34683,I32834,g34688,
    I32837,g34689,I32840,g34690,I32843,g34691,I32846,g34692,g34697,g34698,I32855,g34699,
    g34711,I32868,g34712,I32871,g34713,I32874,g34714,I32878,g34716,I32881,g34717,I32884,
    g34718,I32904,g34736,I32909,g34739,I32921,g34749,I32929,g34755,I32935,g34759,I32938,
    g34760,g34766,I32947,g34767,I32950,g34768,I32953,g34769,I32956,g34770,I32960,g34772,
    I32963,g34773,I32967,g34775,I32970,g34776,I32973,g34777,I32976,g34778,I32982,g34784,
    I32985,g34785,I32988,g34786,I32991,g34787,I32994,I32997,g34789,I33020,g34810,I33024,
    g34812,I33027,g34813,I33030,g34816,I33034,g34820,I33037,g34823,I33041,g34827,I33044,
    g34830,I33047,g34833,I33050,g34836,I33053,I33056,g34840,g34844,g34845,I33064,g34846,
    I33067,g34847,I33070,g34848,I33075,g34851,g34852,I33079,g34855,g34864,I33103,g34877,
    I33106,g34878,I33109,g34879,g34883,I33119,g34893,g34910,I33131,I33134,g34914,I33137,
    I33140,g34916,I33143,I33146,g34918,I33149,I33152,g34920,I33155,I33158,g34922,I33161,
    I33164,g34924,I33167,I33170,g34926,I33173,I33176,g34928,I33179,g34929,I33182,g34930,
    g34932,g34933,g34934,I33189,g34935,g34938,g34939,g34940,g34941,g34942,I33197,g34943,
    g34944,g34945,g34946,g34947,g34949,g34950,g34951,g34952,I33210,g34954,I33214,I33218,
    g34960,I33232,I33235,g34973,g34981,I33246,g34982,I33249,g34983,I33252,g34984,I33255,
    g34985,I33258,g34986,I33261,g34987,I33264,g34988,I33267,g34989,I33270,g34990,I33273,
    g34991,I33276,g34992,I33279,g34993,I33282,g34994,I33285,g34995,I33288,g34996,I33291,
    g34997,g34998,I33297,g35001,I33300,g35002,g7251,g7396,g7469,g7511,g7520,g7685,g7696,
    g7763,g7777,g7804,g7918,g7948,g8234,g8530,g8583,g8643,g8690,g8721,g9217,g9479,g9906,
    g9967,g9968,g10034,g10290,I13862,g10476,g10501,g10528,g10543,g10565,g10588,I13937,
    g10590,g10616,g10619,g10624,g10625,g10626,g10632,g10654,g10655,g10656,g10657,g10665,
    g10674,g10675,g10676,g10677,g10683,g10684,g10704,g10705,g10706,g10707,g10719,g10720,
    g10721,g10724,g10732,g10733,g10736,g10756,g10822,g10823,g10827,g10828,g10829,g10838,
    g10841,g10856,g10869,g10873,g10874,g10878,g10883,g10887,g10890,g10896,g10898,g10902,
    g10917,g10921,g10925,g10934,g10947,g10948,g10966,g10967,g10970,g10998,g10999,g11003,
    g11010,g11016,g11018,g11019,g11023,g11024,g11027,g11028,g11029,g11032,g11035,g11036,
    g11037,g11044,g11045,g11046,g11047,g11083,g11111,g11114,g11115,g11116,g11123,g11126,
    g11127,g11139,g11142,I14198,g11144,g11160,g11163,I14225,g11166,g11178,g11205,g11223,
    g11244,g11366,g11397,g11427,g11449,g11496,g11497,g11546,g11740,g11890,g11893,g11915,
    g11916,g11937,g11939,g11956,g11960,g11967,g11978,g12015,g12027,g12043,g12065,g12099,
    g12135,g12179,g12186,g12219,g12220,g12259,g12284,g12527,g12641,g12687,g12692,g12730,
    g12735,g12761,g12762,g12794,g12795,g12812,g12817,g12920,g12924,g12931,g12939,g12953,
    g12979,g13019,g13020,g13025,g13029,g13030,g13035,g13038,g13042,g13046,g13047,g13048,
    g13059,g13060,g13063,g13080,g13081,g13156,g13221,g13247,g13252,g13265,g13277,g13282,
    g13287,g13290,g13294,g13299,g13306,g13313,g13319,g13320,g13321,g13324,g13333,g13345,
    g13349,g13383,g13384,g13393,g13411,g13415,g13436,g13461,g13473,g13491,g13492,g13493,
    g13497,g13507,g13508,g13509,g13523,g13524,g13525,g13541,g13542,g13564,g13566,g13567,
    g13604,g13632,g13633,g13656,g13671,g13697,g13737,g13738,I16111,g13771,g13778,I16129,
    g13805,g13807,g13808,I16143,g13830,g13832,g13833,g13853,g13887,g13912,g13942,g13974,
    g13998,g14028,g14035,g14061,g14097,g14126,g14148,g14168,g14180,g14185,g14190,g14193,
    g14202,g14206,g14207,g14210,g14216,g14218,g14220,g14221,g14222,g14233,g14256,g14257,
    g14261,g14295,g14296,g14316,g14438,I16618,g14496,g14506,I16646,g14528,g14537,I16671,
    g14555,g14565,g14566,g14567,I16695,g14581,g14585,g14586,g14587,g14588,g14589,I16721,
    g14608,g14610,g14612,g14613,g14614,g14615,g14641,g14643,g14644,g14654,g14680,g14681,
    g14708,g14719,g14791,g14831,g14832,g14874,g14875,g14913,g15075,g15076,g15077,g15078,
    g15079,g15080,g15081,g15082,g15083,g15084,g15103,g15104,g15105,g15107,g15108,g15109,
    g15110,g15111,g15112,g15113,g15114,g15115,g15116,g15117,g15118,g15119,g15507,g15567,
    g15574,g15589,g15590,g15611,g15612,g15613,g15631,g15632,g15633,g15650,g15651,g15652,
    g15653,g15654,g15672,g15673,g15678,g15679,g15693,g15694,g15699,g15700,g15701,g15703,
    g15704,g15706,g15707,g15711,g15712,g15716,g15722,g15738,g15745,g15749,g15757,g15779,
    g15783,g15784,g15785,g15786,g15793,g15794,g15795,g15796,g15797,g15804,g15805,g15807,
    g15808,g15809,g15810,g15812,g15813,g15814,g15815,g15817,g15818,g15819,g15820,g15821,
    g15822,g15823,g15836,g15837,g15838,g15839,g15840,g15841,g15847,g15848,g15849,g15850,
    g15851,g15852,g15856,g15857,g15858,g15859,g15860,g15861,g15863,g15870,g15871,g15872,
    g15873,g15874,g15875,g15876,g15880,g15881,g15882,g15883,g15884,g15902,g15903,g15911,
    g15912,g15913,g15914,g15936,g15937,g15966,g15967,g15978,g15995,g16023,g16025,g16026,
    g16047,g16098,g16122,g16125,g16126,g16128,g16160,g16161,g16163,g16176,g16177,g16178,
    g16179,g16184,g16185,g16190,g16191,g16192,g16193,I17529,g16194,g16199,g16202,g16203,
    g16204,I17542,g16205,g16207,g16208,g16211,g16212,I17552,g16213,g16221,g16222,g16224,
    g16233,I17575,g16234,g16243,I17585,g16244,g16245,g16279,I17606,g16283,g16303,g16324,
    g16422,g16427,g16474,g16483,g16484,g16485,I17692,g16486,g16513,g16516,g16517,g16518,
    g16519,g16520,g16531,g16532,g16534,g16535,g16536,g16537,g16538,I17741,g16539,g16590,
    g16591,g16592,g16593,g16595,g16596,g16597,g16598,g16599,g16610,g16611,g16612,g16613,
    g16614,g16616,g16617,g16618,g16619,g16621,g16633,g16634,g16635,g16636,g16637,g16638,
    g16639,g16641,g16642,g16653,g16662,g16666,g16667,g16668,g16669,g16670,g16671,g16672,
    g16673,g16674,g16690,g16699,g16700,g16701,g16702,g16703,g16704,g16705,g16706,g16707,
    g16729,g16730,g16731,g16732,g16733,g16734,g16735,g16736,g16737,g16751,g16758,g16759,
    g16760,g16761,g16762,g16763,g16764,g16765,g16766,g16801,g16802,g16803,g16804,g16805,
    g16806,g16807,g16808,g16840,g16841,g16842,g16843,g16844,g16845,g16846,g16855,g16868,
    g16869,g16870,g16871,g16884,g16885,g16896,g16929,g16930,g16957,g16965,g16986,g17057,
    g17091,g17119,g17123,g17133,g17134,g17138,g17139,g17140,g17145,g17146,g17149,g17150,
    g17151,g17152,g17153,g17156,g17176,g17177,g17179,g17181,g17182,g17191,g17192,g17193,
    g17199,g17292,g17307,g17317,g17321,g17365,g17391,g17401,g17405,g17418,g17424,g17469,
    g17480,g17506,g17574,g17601,I18568,g17613,g17617,g17636,g17643,I18620,g17653,g17654,
    g17655,g17671,g17682,I18671,g17690,g17692,g17693,g17719,I18713,g17724,I18716,g17725,
    g17726,I18740,g17747,g17752,g17753,I18762,g17766,I18765,g17767,g17768,g17769,g17770,
    g17771,I18782,g17780,I18785,g17781,g17783,g17784,g17785,g17786,I18803,g17793,g17809,
    g17810,I18819,g17817,g18103,g18104,g18105,g18106,g18107,g18108,g18109,g18110,g18111,
    g18112,g18113,g18114,g18115,g18116,g18117,g18118,g18119,g18120,g18121,g18122,g18123,
    g18124,g18125,g18126,g18127,g18128,g18129,g18130,g18131,g18132,g18133,g18134,g18135,
    g18136,g18137,g18138,g18139,g18140,g18141,g18142,g18143,g18144,g18145,g18146,g18147,
    g18148,g18149,g18150,g18151,g18152,g18153,g18154,g18155,g18156,g18157,g18158,g18159,
    g18160,g18161,g18162,g18163,g18164,g18165,g18166,g18167,g18168,g18169,g18170,g18171,
    g18172,g18173,g18174,g18175,g18176,g18177,g18178,g18179,g18180,g18181,g18182,g18183,
    g18184,g18185,g18186,g18187,g18188,g18189,g18190,g18191,g18192,g18193,g18194,g18195,
    g18196,g18197,g18198,g18199,g18201,g18202,g18203,g18204,g18205,g18206,g18207,g18208,
    g18209,g18210,g18211,g18212,g18213,g18214,g18215,g18216,g18217,g18218,g18219,g18220,
    g18221,g18222,g18223,g18224,g18225,g18226,g18227,g18228,g18229,g18230,g18231,g18232,
    g18233,g18234,g18235,g18236,g18237,g18238,g18239,g18240,g18241,g18242,g18243,g18244,
    g18245,g18246,g18247,g18248,g18249,g18250,g18251,g18252,g18253,g18254,g18255,g18256,
    g18257,g18258,g18259,g18260,g18261,g18262,g18263,g18264,g18265,g18266,g18267,g18268,
    g18269,g18270,g18271,g18272,g18273,g18274,g18275,g18276,g18277,g18278,g18279,g18280,
    g18281,g18282,g18283,g18284,g18285,g18286,g18287,g18288,g18289,g18290,g18291,g18292,
    g18293,g18294,g18295,g18296,g18297,g18298,g18299,g18300,g18301,g18302,g18303,g18304,
    g18305,g18306,g18307,g18308,g18309,g18310,g18311,g18312,g18313,g18314,g18315,g18316,
    g18317,g18318,g18319,g18320,g18321,g18322,g18323,g18324,g18325,g18326,g18327,g18328,
    g18329,g18330,g18331,g18332,g18333,g18334,g18335,g18336,g18337,g18338,g18339,g18340,
    g18341,g18342,g18343,g18344,g18345,g18346,g18347,g18348,g18349,g18350,g18351,g18352,
    g18353,g18354,g18355,g18356,g18357,g18358,g18359,g18360,g18361,g18362,g18363,g18364,
    g18365,g18366,g18367,g18368,g18369,g18370,g18371,g18372,g18373,g18374,g18375,g18376,
    g18377,g18378,g18379,g18380,g18381,g18382,g18383,g18384,g18385,g18386,g18387,g18388,
    g18389,g18390,g18391,g18392,g18393,g18394,g18395,g18396,g18397,g18398,g18399,g18400,
    g18401,g18402,g18403,g18404,g18405,g18406,g18407,g18408,g18409,g18410,g18411,g18412,
    g18413,g18414,g18415,g18416,g18417,g18418,g18419,g18420,g18423,g18424,g18425,g18426,
    g18427,g18428,g18429,g18430,g18431,g18432,g18433,g18434,g18435,g18436,g18437,g18438,
    g18439,g18440,g18441,g18442,g18443,g18444,g18445,g18446,g18447,g18448,g18449,g18450,
    g18451,g18452,g18453,g18454,g18455,g18456,g18457,g18458,g18459,g18460,g18461,g18462,
    g18463,g18464,g18465,g18466,g18467,g18468,g18469,g18470,g18471,g18472,g18473,g18474,
    g18475,g18476,g18477,g18478,g18479,g18480,g18481,g18482,g18483,g18484,g18485,g18486,
    g18487,g18488,g18489,g18490,g18491,g18492,g18493,g18494,g18495,g18496,g18497,g18498,
    g18499,g18500,g18501,g18502,g18503,g18504,g18505,g18506,g18507,g18508,g18509,g18510,
    g18511,g18512,g18513,g18514,g18515,g18516,g18517,g18518,g18519,g18520,g18521,g18522,
    g18523,g18524,g18525,g18526,g18529,g18530,g18531,g18532,g18533,g18534,g18535,g18536,
    g18537,g18538,g18539,g18540,g18541,g18542,g18543,g18544,g18545,g18546,g18547,g18548,
    g18549,g18550,g18551,g18552,g18553,g18554,g18555,g18556,g18557,g18558,g18559,g18560,
    g18561,g18563,g18564,g18565,g18566,g18567,g18568,g18569,g18570,g18571,g18572,g18573,
    g18574,g18575,g18576,g18577,g18578,g18579,g18580,g18581,g18582,g18583,g18584,g18585,
    g18586,g18587,g18588,g18589,g18590,g18591,g18592,g18593,g18594,g18595,g18596,g18597,
    g18598,g18599,g18600,g18601,g18602,g18603,g18604,g18605,g18606,g18607,g18608,g18609,
    g18610,g18611,g18612,g18613,g18614,g18615,g18616,g18617,g18618,g18619,g18620,g18621,
    g18622,g18623,g18624,g18625,g18626,g18627,g18628,g18629,g18630,g18631,g18632,g18633,
    g18634,g18635,g18636,g18637,g18638,g18639,g18640,g18641,g18642,g18643,g18644,g18645,
    g18646,g18647,g18648,g18649,g18650,g18651,g18652,g18653,g18654,g18655,g18656,g18657,
    g18658,g18659,g18662,g18663,g18664,g18665,g18666,g18667,g18668,g18669,g18670,g18671,
    g18672,g18673,g18674,g18675,g18676,g18677,g18678,g18679,g18680,g18681,g18682,g18683,
    g18684,g18685,g18686,g18687,g18688,g18689,g18690,g18691,g18692,g18693,g18694,g18695,
    g18696,g18697,g18698,g18699,g18700,g18701,g18702,g18703,g18704,g18705,g18706,g18707,
    g18708,g18709,g18710,g18711,g18712,g18713,g18714,g18715,g18716,g18717,g18718,g18719,
    g18720,g18721,g18722,g18723,g18724,g18725,g18726,g18727,g18728,g18729,g18730,g18731,
    g18732,g18733,g18734,g18735,g18736,g18737,g18738,g18739,g18740,g18741,g18742,g18743,
    g18744,g18745,g18746,g18747,g18748,g18749,g18750,g18751,g18752,g18753,g18754,g18755,
    g18756,g18757,g18758,g18759,g18760,g18761,g18762,g18763,g18764,g18765,g18766,g18767,
    g18768,g18769,g18770,g18771,g18772,g18773,g18774,g18775,g18776,g18777,g18778,g18779,
    g18780,g18781,g18782,g18783,g18784,g18785,g18786,g18787,g18788,g18789,g18790,g18791,
    g18792,g18793,g18794,g18795,g18796,g18797,g18798,g18799,g18800,g18801,g18802,g18803,
    g18804,g18805,g18806,g18807,g18808,g18809,g18810,g18811,g18812,g18813,g18814,g18815,
    g18816,g18817,g18818,g18819,g18820,g18821,g18822,g18823,g18824,g18825,g18826,g18890,
    g18893,g18906,g18909,g18910,g18933,g18934,g18935,g18943,g18949,g18950,g18951,g18974,
    g18981,g18982,g18987,g18992,g18993,g19062,g19069,g19139,g19145,g19206,g19207,g19266,
    g19275,g19333,g19350,g19354,g19372,g19383,g19384,g19393,g19461,g19462,g19487,g19500,
    g19516,g19521,g19536,g19540,g19545,g19556,g19560,g19564,g19568,g19571,g19578,g19581,
    g19585,g19588,g19594,g19596,g19601,g19610,g19613,g19631,g19637,g19651,g19655,g19656,
    g19660,g19661,g19671,g19674,g19680,g19681,g19684,g19691,g19692,g19693,g19715,g19716,
    g19717,g19735,g19736,g19740,g19746,g19749,g19752,g19756,g19767,g19768,g19784,g19788,
    g19791,g19855,g19911,g19914,g19948,g20056,g20069,g20084,g20093,g20094,g20095,g20108,
    g20109,g20112,g20131,g20135,g20152,g20162,g20165,g20171,g20174,g20188,g20193,g20203,
    g20215,g20218,g20375,g20559,g20581,g20602,g20628,g20658,g20682,g20739,g20751,g20875,
    g20887,g20977,g21012,g21024,g21066,g21067,g21163,g21188,g21251,g21276,g21285,g21296,
    g21298,g21302,g21303,g21332,g21333,g21347,g21348,g21361,g21378,g21382,g21394,g21404,
    g21405,g21419,g21420,g21452,g21453,g21464,g21465,g21512,g21513,g21557,g21558,g21559,
    g21605,g21606,g21699,g21700,g21701,g21702,g21703,g21704,g21705,g21706,g21707,g21708,
    g21709,g21710,g21711,g21712,g21713,g21714,g21715,g21716,g21717,g21718,g21719,g21720,
    g21721,g21728,g21729,g21730,g21731,g21732,g21733,g21734,g21735,g21736,g21737,g21738,
    g21739,g21740,g21741,g21742,g21743,g21744,g21745,g21746,g21747,g21748,g21749,g21750,
    g21751,g21752,g21753,g21754,g21755,g21756,g21757,g21758,g21759,g21760,g21761,g21762,
    g21763,g21764,g21765,g21766,g21767,g21768,g21769,g21770,g21771,g21772,g21773,g21774,
    g21775,g21776,g21777,g21778,g21779,g21780,g21781,g21782,g21783,g21784,g21785,g21786,
    g21787,g21788,g21789,g21790,g21791,g21792,g21793,g21794,g21795,g21796,g21797,g21798,
    g21799,g21800,g21801,g21802,g21803,g21804,g21805,g21806,g21807,g21808,g21809,g21810,
    g21811,g21812,g21813,g21814,g21815,g21816,g21817,g21818,g21819,g21820,g21821,g21822,
    g21823,g21824,g21825,g21826,g21827,g21828,g21829,g21830,g21831,g21832,g21833,g21834,
    g21835,g21836,g21837,g21838,g21839,g21840,g21841,g21842,g21843,g21844,g21845,g21846,
    g21847,g21848,g21849,g21850,g21851,g21852,g21853,g21854,g21855,g21856,g21857,g21858,
    g21859,g21860,g21861,g21862,g21863,g21864,g21865,g21866,g21867,g21868,g21869,g21870,
    g21871,g21872,g21873,g21874,g21875,g21876,g21877,g21878,g21879,g21880,g21881,g21882,
    g21883,g21884,g21885,g21886,g21887,g21888,g21889,g21890,g21906,g21907,g21908,g21909,
    g21910,g21911,g21912,g21913,g21914,g21915,g21916,g21917,g21918,g21919,g21920,g21921,
    g21922,g21923,g21924,g21925,g21926,g21927,g21928,g21929,g21930,g21931,g21932,g21933,
    g21934,g21935,g21936,g21937,g21938,g21939,g21940,g21941,g21942,g21943,g21944,g21945,
    g21946,g21947,g21948,g21949,g21950,g21951,g21952,g21953,g21954,g21955,g21956,g21957,
    g21958,g21959,g21960,g21961,g21962,g21963,g21964,g21965,g21966,g21967,g21968,g21969,
    g21970,g21971,g21972,g21973,g21974,g21975,g21976,g21977,g21978,g21979,g21980,g21981,
    g21982,g21983,g21984,g21985,g21986,g21987,g21988,g21989,g21990,g21991,g21992,g21993,
    g21994,g21995,g21996,g21997,g21998,g21999,g22000,g22001,g22002,g22003,g22004,g22005,
    g22006,g22007,g22008,g22009,g22010,g22011,g22012,g22013,g22014,g22015,g22016,g22017,
    g22018,g22019,g22020,g22021,g22022,g22023,g22024,g22025,g22026,g22027,g22028,g22029,
    g22030,g22031,g22032,g22033,g22034,g22035,g22036,g22037,g22038,g22039,g22040,g22041,
    g22042,g22043,g22044,g22045,g22046,g22047,g22048,g22049,g22050,g22051,g22052,g22053,
    g22054,g22055,g22056,g22057,g22058,g22059,g22060,g22061,g22062,g22063,g22064,g22065,
    g22066,g22067,g22068,g22069,g22070,g22071,g22072,g22073,g22074,g22075,g22076,g22077,
    g22078,g22079,g22080,g22081,g22082,g22083,g22084,g22085,g22086,g22087,g22088,g22089,
    g22090,g22091,g22092,g22093,g22094,g22095,g22096,g22097,g22098,g22099,g22100,g22101,
    g22102,g22103,g22104,g22105,g22106,g22107,g22108,g22109,g22110,g22111,g22112,g22113,
    g22114,g22115,g22116,g22117,g22118,g22119,g22120,g22121,g22122,g22123,g22124,g22125,
    g22126,g22127,g22128,g22129,g22130,g22131,g22132,g22133,g22134,g22135,g22142,g22143,
    g22145,g22149,g22157,g22158,g22160,g22161,g22165,g22172,g22191,g22193,g22208,g22209,
    g22216,g22218,g22219,g22298,g22299,g22307,g22308,g22309,g22310,g22316,g22329,g22340,
    g22342,g22369,g22384,g22417,g22432,g22457,g22472,g22489,g22498,g22515,g22518,g22525,
    g22534,g22538,g22588,g22589,g22590,g22622,g22623,g22624,g22632,g22633,g22637,g22665,
    g22670,g22680,g22685,g22686,g22689,g22710,g22717,g22720,g22752,g22760,g22762,g22831,
    g22834,g22835,g22843,g22846,g22848,g22849,g22851,g22859,g22861,g22862,g22863,g22871,
    g22873,g22876,g22899,g22900,g22920,g22937,g22938,g22939,g22942,g22982,g22990,g22991,
    g22992,g23006,g23007,g23008,g23009,g23023,g23025,g23050,g23056,g23062,g23076,g23083,
    g23103,g23104,g23121,g23130,g23131,g23148,g23151,g23165,g23166,g23187,g23188,g23201,
    g23218,g23220,g23229,g23254,g23265,g23280,g23292,g23293,g23314,g23348,g23349,g23372,
    g23373,g23381,g23386,g23387,g23389,g23392,g23396,g23397,g23401,g23404,g23407,g23412,
    g23415,g23416,g23424,g23436,g23439,g23451,g23471,g23474,g23475,g23484,g23497,g23498,
    g23513,g23514,g23531,g23532,g23533,g23540,g23551,g23553,g23554,g23564,g23572,g23577,
    g23581,g23599,g23606,g23618,g23619,g23639,g23646,g23657,g23658,g23675,g23682,g23690,
    g23691,g23708,g23724,g23725,g23742,g23754,g23755,g23774,g23775,g23779,g23799,g23801,
    g23802,g23811,g23828,g23836,g23837,g23854,g23855,g23856,g23857,g23872,g23873,g23884,
    g23885,g23900,g23901,g23917,g23919,g23920,g23921,g23957,g23958,g23990,g23991,g23996,
    g23998,g24001,g24002,g24004,g24008,g24009,g24011,g24012,g24014,g24015,g24016,g24139,
    g24140,g24141,g24142,g24143,g24144,g24186,g24187,g24188,g24189,g24190,g24191,g24192,
    g24193,g24194,g24195,g24196,g24197,g24198,g24199,g24217,g24218,g24219,g24220,g24221,
    g24222,g24223,g24224,g24225,g24226,g24227,g24228,g24229,g24230,g24283,g24284,g24285,
    g24286,g24287,g24288,g24289,g24290,g24291,g24292,g24293,g24294,g24295,g24296,g24297,
    g24298,g24299,g24300,g24301,g24302,g24303,g24304,g24305,g24306,g24307,g24308,g24309,
    g24310,g24311,g24312,g24313,g24314,g24315,g24316,g24317,g24318,g24319,g24320,g24321,
    g24322,g24323,g24324,g24325,g24326,g24327,g24328,g24329,g24330,g24331,g24332,g24333,
    g24378,g24387,g24392,g24393,g24395,g24399,g24400,g24402,g24403,g24406,g24408,g24409,
    g24410,g24411,g24415,g24416,g24420,g24421,g24422,g24423,g24427,g24436,g24450,g24451,
    g24464,g24465,g24467,g24475,g24476,g24482,g24484,g24485,g24488,g24491,g24495,g24498,
    g24499,g24501,g24502,g24503,g24504,g24507,g24523,g24532,g24536,g24537,g24541,g24545,
    g24546,g24549,g24550,g24551,g24552,g24553,g24554,g24555,g24556,g24558,g24559,g24564,
    g24569,g24572,g24573,g24581,g24582,g24588,g24589,g24590,g24600,g24602,g24606,g24607,
    g24608,g24618,g24622,g24624,g24627,g24628,g24629,g24630,g24634,g24635,g24637,g24638,
    g24639,g24640,g24642,g24643,g24644,g24645,g24646,g24647,g24649,g24650,g24651,g24654,
    g24656,g24657,g24658,g24659,g24660,g24663,g24664,g24666,g24668,g24669,g24670,g24671,
    g24672,g24673,g24674,g24675,g24676,g24679,g24680,g24681,g24682,g24684,g24686,g24687,
    g24688,g24698,g24700,g24702,g24703,g24704,g24706,g24707,g24708,g24709,g24710,g24712,
    g24713,g24714,g24716,g24717,g24719,g24721,g24722,g24723,g24724,g24725,g24726,g24727,
    g24728,g24729,g24730,g24731,g24743,g24745,g24747,g24748,g24749,g24750,g24754,g24755,
    g24757,g24758,g24761,g24762,g24763,g24764,g24765,g24769,g24771,g24772,g24773,g24774,
    g24775,g24777,g24785,g24786,g24788,g24790,g24794,g24796,g24797,g24803,g24812,g24817,
    g24820,I24003,g24822,g24835,I24015,g24843,I24018,g24846,g24849,I24027,g24855,I24030,
    g24858,I24033,g24861,g24864,g24865,g24872,I24048,g24881,I24051,g24884,I24054,g24887,
    g24892,I24064,g24897,I24067,g24900,g24903,g24904,I24075,g24908,g24912,g24913,g24914,
    g24915,g24921,g24922,g24923,g24929,g24930,g24931,g24939,g24940,g24941,g24945,g24949,
    g24961,g24962,g24967,g24977,g24983,g24984,g24997,g24998,g25012,g25014,g25026,g25030,
    g25031,g25033,g25040,g25041,g25042,g25043,g25045,g25050,g25054,g25056,g25057,g25058,
    g25059,g25061,g25063,g25067,g25068,g25069,g25071,g25076,g25077,g25078,g25079,g25084,
    g25085,g25086,g25087,g25088,g25089,g25091,g25093,g25094,g25095,g25096,g25102,g25103,
    g25104,g25105,g25106,g25107,g25108,g25110,g25112,g25113,g25122,g25123,g25124,g25125,
    g25126,g25127,g25128,g25129,g25130,g25132,g25142,g25143,g25147,g25148,g25149,g25150,
    g25151,g25152,g25159,g25163,g25164,g25165,g25166,g25173,g25178,g25179,g25181,g25187,
    g25192,g25201,g25207,g25217,g25223,g25229,g25238,g25285,I24482,g25290,g25323,I24505,
    g25328,I24508,g25331,g25357,g25366,g25367,g25368,I24524,g25371,I24527,g25374,I24530,
    g25377,g25408,I24546,g25411,I24549,g25414,I24552,g25417,I24555,g25420,g25448,g25449,
    g25450,I24576,g25453,I24579,g25456,I24582,g25459,I24585,g25462,g25466,g25479,I24597,
    g25482,I24600,g25485,I24603,g25488,g25491,g25502,g25503,I24616,g25507,I24619,g25510,
    I24625,g25518,g25522,g25526,g25530,g25536,g25543,g25551,g25559,g25565,I24674,I24675,
    g25567,I24679,I24680,g25568,I24684,I24685,g25569,I24689,I24690,g25570,I24694,I24695,
    g25571,I24699,I24700,g25572,I24704,I24705,g25573,I24709,I24710,g25574,g25578,g25579,
    g25580,g25581,g25765,g25768,g25772,g25775,g25780,g25782,g25787,g25788,g25801,g25802,
    g25803,g25804,g25814,g25815,g25816,g25817,g25818,g25831,g25832,g25833,g25848,g25850,
    g25852,g25865,g25866,g25870,g25871,g25872,g25873,g25874,g25875,g25876,g25879,g25880,
    g25881,g25883,g25884,g25900,g25901,g25902,g25904,g25905,g25907,g25908,g25909,g25915,
    g25916,g25921,g25922,g25923,g25924,g25925,g25926,g25927,g25928,g25931,g25938,g25939,
    g25946,g25949,g25951,g25955,g25957,g25959,g25961,g25962,g25963,g25964,g25965,g25966,
    g25967,g25968,g25969,g25970,g25971,g25972,g25973,g25975,g25976,g25977,g25978,g25979,
    g25980,g25981,g25982,g25983,g25986,g25987,g25988,g25989,g25990,g25991,g25992,g25993,
    g26019,g26020,g26021,g26022,g26023,g26024,g26048,g26049,g26050,g26051,g26077,g26078,
    g26079,g26084,g26085,g26086,g26087,g26088,g26090,g26091,g26092,g26094,g26095,g26096,
    g26097,g26100,g26101,g26102,g26103,g26104,g26119,g26120,g26121,g26122,g26123,g26124,
    g26125,g26126,g26127,g26128,g26129,g26130,g26145,g26146,g26147,g26148,g26153,g26154,
    g26155,g26156,g26157,g26158,g26159,g26160,g26161,g26165,g26166,g26171,g26176,g26177,
    g26178,g26179,g26180,g26181,g26182,g26186,g26190,g26195,g26200,g26203,g26204,g26205,
    g26206,g26207,g26213,g26218,g26223,g26226,g26229,g26230,g26231,g26232,g26233,g26234,
    g26236,g26241,g26244,g26249,g26250,g26251,g26252,g26253,g26254,g26257,g26258,g26259,
    g26261,g26264,g26270,g26271,g26272,g26273,g26274,g26275,g26276,g26277,g26279,g26280,
    g26281,g26285,g26286,g26287,g26288,g26289,g26290,g26291,g26292,g26294,g26295,g26300,
    g26301,g26302,g26303,g26304,g26306,g26307,g26308,g26310,g26311,g26312,g26313,g26323,
    g26324,g26325,g26336,g26339,g26341,g26345,g26347,g26350,g26351,g26356,g26357,g26358,
    g26360,g26362,g26378,g26379,g26380,g26381,g26387,g26388,g26389,g26390,g26391,g26393,
    g26394,g26395,g26397,g26398,g26399,g26423,g26484,g26485,g26486,g26487,g26511,g26513,
    g26514,g26516,g26517,g26541,g26542,g26543,g26544,g26547,g26571,g26572,g26602,g26604,
    g26606,g26610,g26611,g26612,g26613,g26629,g26630,g26633,g26635,g26650,g26651,g26652,
    g26670,g26671,g26684,g26689,g26711,g26712,g26713,g26719,g26749,g26750,g26753,g26778,
    g26779,g26780,g26783,g26799,g26808,g26815,g26819,g26821,g26822,g26823,g26826,g26828,
    g26829,g26833,g26838,g26839,g26842,g26844,g26845,g26846,g26847,g26848,g26849,g26852,
    g26853,g26854,g26855,g26857,g26858,g26861,g26863,g26864,g26871,g26977,g26994,g27020,
    g27025,g27028,g27029,g27030,g27032,g27033,g27034,g27035,g27036,g27039,g27040,g27041,
    g27042,g27043,g27044,g27045,g27050,g27057,g27058,g27073,g27083,g27085,g27086,g27087,
    g27090,g27094,g27095,g27096,g27097,g27098,g27099,g27103,g27104,g27105,g27106,g27107,
    g27113,g27114,g27115,g27116,g27117,g27118,g27119,g27120,g27121,g27127,g27128,g27129,
    g27130,g27131,g27132,g27134,g27136,g27137,g27138,g27139,g27140,g27145,g27146,g27148,
    g27149,g27151,g27153,g27154,g27158,g27160,g27161,g27162,g27177,g27178,g27180,g27181,
    g27183,g27184,g27185,g27186,g27201,g27202,g27203,g27204,g27206,g27207,g27208,g27209,
    g27210,g27211,g27212,g27213,g27214,g27215,g27216,g27217,g27218,g27219,g27220,g27221,
    g27222,g27227,g27228,g27229,g27230,g27234,g27235,g27246,g27247,g27249,g27251,g27252,
    g27254,g27255,g27256,g27259,g27260,g27262,g27263,g27264,g27265,g27266,g27267,g27268,
    g27269,g27270,g27272,g27275,g27276,g27277,g27280,g27281,g27284,g27285,g27286,g27287,
    g27288,g27291,g27292,g27293,g27294,g27298,g27299,g27300,g27301,g27302,g27303,g27304,
    g27305,g27309,g27310,g27311,g27312,g27313,g27314,g27315,g27316,g27323,g27324,g27325,
    g27326,g27327,g27328,g27329,g27330,g27331,g27332,g27333,g27334,g27335,g27336,g27339,
    g27340,g27341,g27342,g27346,g27347,g27348,g27350,g27351,g27357,g27358,g27359,g27360,
    g27361,g27362,g27363,g27369,g27370,g27371,g27372,g27373,g27374,g27375,g27376,g27378,
    g27384,g27385,g27386,g27387,g27388,g27389,g27390,g27391,g27392,g27393,g27395,g27404,
    g27406,g27407,g27408,g27409,g27410,g27411,g27412,g27413,g27414,g27416,g27421,g27427,
    g27428,g27430,g27432,g27433,g27434,g27435,g27436,g27437,g27439,g27440,g27445,g27451,
    g27452,g27454,g27455,g27457,g27459,g27460,g27461,g27462,g27467,g27469,g27474,g27480,
    g27481,g27482,g27483,g27485,g27486,g27488,g27490,g27491,g27493,g27494,g27500,g27501,
    g27502,g27503,g27504,g27505,g27507,g27508,g27510,g27517,g27518,g27519,g27520,g27521,
    g27522,g27523,g27525,g27526,g27534,g27535,g27536,g27537,g27538,g27539,g27540,g27541,
    g27545,g27546,g27547,g27548,g27549,g27553,g27557,g27558,g27559,g27560,g27564,g27568,
    g27588,g27594,g27595,g27598,g27599,g27600,g27601,g27602,g27612,g27614,g27615,g27616,
    g27617,g27627,g27628,g27633,g27634,g27635,g27645,g27646,g27648,g27649,g27650,g27651,
    g27653,g27658,g27660,g27661,g27664,g27665,g27666,g27667,g27668,g27669,g27673,g27674,
    g27676,g27677,g27678,g27682,g27683,g27684,g27685,g27686,g27690,g27691,g27692,g27696,
    g27697,g27699,g27700,g27710,g27711,g27714,g27723,g27724,g27727,g27759,g27762,g27765,
    g27817,g27820,g27821,g27822,g27932,g27957,g27958,g27959,g27962,g27963,g27964,g27965,
    g27968,g27981,g27988,g27992,g27995,g27997,g27999,g28010,g28020,I26530,I26531,g28035,
    g28107,g28108,g28110,g28111,g28112,g28113,g28114,g28115,g28116,g28117,g28124,g28125,
    g28130,g28133,g28136,g28139,g28141,g28143,g28144,g28148,g28150,g28151,g28152,g28153,
    g28154,g28158,g28159,g28160,g28164,g28165,g28171,g28178,g28182,g28183,g28185,g28192,
    g28193,g28197,g28198,g28199,g28200,g28201,g28202,g28204,g28205,g28210,g28213,g28214,
    g28215,g28217,g28218,g28219,g28223,g28224,g28225,g28226,g28227,g28228,g28229,g28231,
    g28232,g28233,g28234,g28235,g28236,g28237,g28238,g28239,g28240,g28242,g28243,g28244,
    g28245,g28246,g28247,g28248,g28249,g28251,g28252,g28253,g28254,g28255,g28256,g28257,
    g28258,g28260,g28261,g28263,g28264,g28265,g28266,g28267,g28268,g28269,g28272,g28273,
    g28280,g28281,g28282,g28283,g28284,g28285,g28289,g28290,g28291,g28292,g28293,g28299,
    g28300,g28301,g28302,g28303,g28304,g28311,g28312,g28313,g28314,g28315,g28318,g28324,
    g28327,g28330,g28333,g28339,g28341,g28343,g28346,g28352,g28360,g28415,g28426,g28427,
    g28439,g28440,g28442,g28451,g28453,g28454,g28455,g28456,I26948,g28458,g28466,g28467,
    I26960,g28471,g28477,g28478,I26972,g28484,g28488,g28489,g28494,g28495,g28499,g28523,
    g28524,g28528,g28530,g28531,g28532,g28535,g28537,g28539,g28541,g28542,g28543,g28547,
    g28550,g28553,g28554,g28555,g28556,g28557,g28558,g28563,g28567,g28569,g28570,g28571,
    g28572,g28573,g28583,g28585,g28586,g28587,g28588,g28597,g28599,g28601,g28602,g28612,
    g28616,g28617,g28624,g28626,g28627,g28630,g28637,g28638,g28639,g28642,g28645,g28652,
    g28653,g28654,g28655,g28657,g28658,g28660,g28663,g28666,g28672,g28673,g28674,g28676,
    g28677,g28679,g28683,g28686,g28689,g28692,g28694,g28695,g28697,g28703,g28706,g28710,
    g28712,g28714,g28722,g28725,g28739,g28761,g28768,g28789,g28799,g28812,g28813,g28833,
    g28846,g28880,g28889,g28919,g28924,g28939,g28959,g28970,I27349,g28982,g28991,g28998,
    I27364,g29008,g29029,I27381,g29036,I27409,g29073,I27429,g29110,g29178,g29182,g29188,
    g29192,g29199,I27503,I27504,g29201,I27508,I27509,g29202,I27513,I27514,g29203,I27518,
    I27519,g29204,I27523,I27524,g29205,I27528,I27529,g29206,I27533,I27534,g29207,I27538,
    I27539,g29208,g29314,g29315,g29316,g29320,g29321,g29322,g29323,g29324,g29326,g29327,
    g29328,g29329,g29330,g29331,g29332,g29334,g29336,g29337,g29338,g29344,g29345,g29346,
    g29347,g29349,g29350,g29351,g29352,g29354,g29360,g29362,g29363,g29364,g29367,g29369,
    g29375,g29376,g29377,g29378,g29380,g29381,g29382,g29383,g29384,g29475,g29477,g29494,
    g29509,g29510,g29511,g29512,g29513,g29514,g29515,g29516,g29517,g29518,g29519,g29521,
    g29522,g29523,g29524,g29525,g29526,g29527,g29528,g29530,g29531,g29532,g29533,g29534,
    g29535,g29536,g29537,g29538,g29547,g29548,g29549,g29550,g29551,g29552,g29553,g29554,
    g29555,g29563,g29564,g29565,g29566,g29567,g29568,g29569,g29570,g29571,g29572,g29573,
    g29574,g29575,g29576,g29577,g29578,g29579,g29580,g29581,g29582,g29584,g29585,g29586,
    g29587,g29588,g29589,g29590,g29591,g29592,g29593,g29594,g29595,g29596,g29598,g29599,
    g29600,g29601,g29602,g29603,g29604,g29605,g29606,g29607,g29608,g29609,g29610,g29611,
    g29612,g29613,g29614,g29615,g29616,g29617,g29618,g29619,g29620,g29621,g29622,g29623,
    g29624,g29625,g29626,g29627,g29628,g29629,g29630,g29631,g29632,g29633,g29634,g29635,
    g29636,g29637,g29638,g29639,g29640,g29641,g29642,g29644,g29645,g29646,g29647,g29648,
    g29649,g29650,g29651,g29652,g29656,g29661,g29662,g29663,g29664,g29665,g29666,g29667,
    g29668,g29683,g29684,g29685,g29686,g29687,g29688,g29693,g29708,g29709,g29710,g29711,
    g29712,g29718,g29731,g29732,g29733,g29736,g29740,g29742,g29743,g29746,g29747,g29749,
    g29750,g29751,g29752,g29757,g29758,g29759,g29760,g29761,g29762,g29766,g29767,g29769,
    g29770,g29771,g29772,g29773,g29774,g29782,g29783,g29784,g29785,g29787,g29788,g29789,
    g29794,g29795,g29796,g29797,g29798,g29799,g29803,g29804,g29805,g29806,g29807,g29808,
    g29809,g29810,g29834,g29835,g29836,g29837,g29838,g29839,g29840,g29841,g29842,g29843,
    g29844,g29845,g29850,g29851,g29852,g29853,g29854,g29855,g29856,g29857,g29858,g29859,
    g29860,g29861,g29865,g29866,g29867,g29868,g29869,g29870,g29871,g29872,g29874,g29875,
    g29876,g29877,g29880,g29881,g29882,g29883,g29884,g29885,g29887,g29888,g29890,g29891,
    g29894,g29895,g29896,g29899,g29901,g29902,g29907,g29909,g29924,g29926,g29937,g29938,
    g29940,g29943,g29949,g29951,g29952,g29954,g29959,g29962,g29964,g29966,g29968,g29969,
    g29973,g29974,g29975,g29979,g29982,g29984,g29985,g29986,g29987,g29988,g29989,g29990,
    g29991,g29992,g30000,g30001,g30002,g30003,g30004,g30005,g30006,g30007,g30008,g30009,
    g30010,g30011,g30015,g30023,g30024,g30025,g30026,g30027,g30028,g30029,g30030,g30031,
    g30032,g30033,g30034,g30035,g30041,g30042,g30043,g30044,g30045,g30046,g30047,g30048,
    g30049,g30050,g30051,g30056,g30057,g30058,g30059,g30060,g30061,g30062,g30064,g30066,
    g30069,g30070,g30071,g30073,g30075,g30078,g30080,g30082,g30083,g30084,g30086,g30089,
    g30091,g30094,g30095,g30096,g30098,g30099,g30101,g30107,g30108,g30109,g30110,g30111,
    g30112,g30118,g30120,g30121,g30122,g30124,g30125,g30126,g30131,g30133,g30135,g30137,
    g30138,g30139,g30140,g30145,g30149,g30151,g30152,g30153,g30154,g30158,g30161,g30164,
    g30165,g30166,g30167,g30168,g30172,g30173,g30174,g30175,g30177,g30178,g30179,g30180,
    g30181,g30185,g30186,g30187,g30188,g30190,g30191,g30192,g30193,g30194,g30196,g30197,
    g30198,g30199,g30200,g30202,g30203,g30204,g30205,g30207,g30208,g30209,g30210,g30211,
    g30212,g30213,g30215,g30216,g30219,g30220,g30221,g30222,g30223,g30224,g30225,g30226,
    g30227,g30228,g30229,g30230,g30231,g30232,g30233,g30234,g30235,g30236,g30238,g30239,
    g30241,g30242,g30243,g30244,g30245,g30246,g30247,g30248,g30250,g30251,g30253,g30254,
    g30255,g30256,g30257,g30258,g30261,g30263,g30264,g30266,g30267,g30268,g30269,g30272,
    g30274,g30275,g30277,g30278,g30281,g30283,g30284,g30289,g30308,g30315,g30316,g30564,
    g30566,g30576,g30577,g30583,g30589,g30590,g30592,g30594,g30595,g30596,g30598,g30599,
    g30600,g30604,g30607,g30612,g30614,g30670,g30671,g30673,g30730,g30731,g30735,g30825,
    g30914,g30915,g30918,g30919,g30920,g30921,g30925,g30926,g30927,g30930,g30935,g30936,
    g30937,g30982,g31015,g31016,g31017,g31018,g31019,g31021,g31066,g31067,g31069,g31070,
    g31115,g31118,g31120,g31122,g31123,g31124,g31125,g31128,g31129,g31130,g31131,g31132,
    g31139,g31140,g31141,g31142,g31143,g31145,g31146,g31147,g31148,g31149,g31150,g31151,
    g31152,g31153,g31154,g31166,g31167,g31168,g31169,g31170,g31182,g31183,g31184,g31185,
    g31186,g31187,g31188,g31194,g31206,g31207,g31208,g31209,g31210,g31211,g31212,g31218,
    g31219,g31220,g31222,g31223,g31224,g31225,g31226,g31228,g31229,g31230,g31231,g31232,
    g31237,g31238,g31240,g31242,g31252,g31261,g31266,g31270,g31271,g31272,g31273,g31275,
    g31278,g31280,g31281,g31282,g31283,g31285,g31286,g31290,g31292,g31296,g31297,g31298,
    g31299,g31300,g31301,g31305,g31309,g31310,g31312,g31313,g31314,g31321,g31323,g31324,
    g31327,g31374,g31376,g31467,g31470,g31471,g31475,g31477,g31478,g31480,g31481,g31484,
    g31485,g31486,g31488,g31489,g31490,g31492,g31493,g31494,g31495,g31496,g31497,g31499,
    g31500,g31501,g31502,g31503,g31504,g31505,g31508,g31513,g31514,g31516,g31517,g31518,
    g31519,g31520,g31523,g31524,g31525,g31526,g31527,g31528,g31540,g31541,g31542,g31554,
    g31566,g31579,g31654,g31672,g31707,g31710,g31744,g31746,g31750,g31752,g31756,g31758,
    g31759,g31763,g31765,g31769,g31776,g31777,g31778,g31780,g31784,g31786,g31787,g31788,
    g31789,g31790,g31792,g31933,g31934,g31936,g31940,g31941,g31943,g31944,g31948,g31949,
    g31959,g31960,g31961,g31962,g31963,g31966,g31967,g31968,g31969,g31974,g31975,g31976,
    g31977,g31985,g31986,g31987,g31988,g31989,g31990,g31991,g31992,g31993,g31994,g31995,
    g31996,g32008,g32009,g32010,g32011,g32012,g32013,g32014,g32016,g32018,g32019,g32020,
    g32028,g32029,g32030,g32031,g32032,g32034,g32035,g32036,g32039,g32040,g32041,g32042,
    g32043,g32044,g32045,g32046,g32047,g32048,g32049,g32050,g32051,g32052,g32053,g32054,
    g32055,g32056,g32067,g32068,g32069,g32070,g32071,g32082,g32083,g32084,g32085,g32086,
    g32087,g32088,g32089,g32095,g32096,g32097,g32098,g32103,g32104,g32105,g32106,g32107,
    g32108,g32109,g32110,g32111,g32112,g32113,g32114,g32115,g32116,g32119,g32120,g32121,
    g32122,g32126,g32127,g32128,g32129,g32139,g32140,g32141,g32142,g32143,g32145,g32146,
    g32147,g32148,g32149,g32150,g32151,g32152,g32153,g32154,g32156,g32157,g32158,g32159,
    g32160,g32161,g32162,g32163,g32164,g32165,g32166,g32167,g32168,g32169,g32170,g32171,
    g32172,g32173,g32174,g32175,g32176,g32177,g32178,g32179,g32180,g32181,g32182,g32183,
    g32184,g32187,g32188,g32189,g32190,g32191,g32193,g32194,g32195,g32196,g32197,g32198,
    g32199,g32200,g32203,g32204,g32205,g32206,g32207,g32224,g32232,g32234,g32241,g32242,
    g32244,g32246,g32248,g32254,g32255,g32256,g32258,g32260,g32261,g32263,g32265,g32269,
    g32270,g32272,g32273,g32274,g32276,g32278,g32281,g32282,g32283,g32284,g32286,g32287,
    g32290,g32291,g32292,g32293,g32295,g32300,g32301,g32302,g32303,g32304,g32305,g32306,
    g32307,g32308,g32309,g32310,g32311,g32312,g32313,g32314,g32315,g32316,g32317,g32321,
    g32322,g32323,g32324,g32325,g32326,g32327,g32328,g32330,g32331,g32332,g32333,g32334,
    g32335,g32336,g32337,g32338,g32339,g32340,g32341,g32342,g32343,g32345,g32348,g32350,
    g32356,g32369,g32376,g32396,g32397,g32400,g32401,g32402,g32403,g32409,g32410,g32411,
    g32412,g32413,g32414,g32418,g32419,g32420,g32425,g32428,g33071,g33073,g33074,g33081,
    g33082,g33086,g33087,g33091,g33099,g33101,g33102,g33104,g33105,g33106,g33110,g33111,
    g33113,g33114,g33121,g33122,g33124,g33126,g33186,g33233,g33237,g33239,g33241,g33242,
    g33243,g33244,g33245,g33247,g33248,g33249,g33252,g33263,g33264,g33269,g33304,g33305,
    g33311,g33322,g33327,g33328,g33329,g33330,g33331,g33332,g33333,g33334,g33338,g33339,
    g33340,g33341,g33342,g33343,g33344,g33345,g33349,g33350,g33351,g33352,g33353,g33355,
    g33356,g33357,g33358,g33359,g33360,g33361,g33362,g33363,g33364,g33365,g33366,g33367,
    g33368,g33369,g33370,g33371,g33372,g33373,g33374,g33376,g33379,g33381,g33392,g33399,
    g33400,g33401,g33402,g33403,g33404,g33405,g33406,g33407,g33408,g33409,g33410,g33411,
    g33412,g33414,g33415,g33416,g33417,g33418,g33420,g33421,g33422,g33423,g33425,g33428,
    g33429,g33431,g33433,g33434,g33440,g33441,g33446,g33450,I31001,I31002,g33461,I31006,
    I31007,g33462,I31011,I31012,g33463,I31016,I31017,g33464,I31021,I31022,g33465,I31026,
    I31027,g33466,I31031,I31032,g33467,I31036,I31037,g33468,I31041,I31042,g33469,I31046,
    I31047,g33470,I31051,I31052,g33471,I31056,I31057,g33472,I31061,I31062,g33473,I31066,
    I31067,g33474,I31071,I31072,g33475,I31076,I31077,g33476,I31081,I31082,g33477,I31086,
    I31087,g33478,I31091,I31092,g33479,I31096,I31097,g33480,I31101,I31102,g33481,I31106,
    I31107,g33482,I31111,I31112,g33483,I31116,I31117,g33484,I31121,I31122,g33485,I31126,
    I31127,g33486,I31131,I31132,g33487,I31136,I31137,g33488,I31141,I31142,g33489,I31146,
    I31147,g33490,I31151,I31152,g33491,I31156,I31157,g33492,I31161,I31162,g33493,I31166,
    I31167,g33494,I31171,I31172,g33495,I31176,I31177,g33496,I31181,I31182,g33497,I31186,
    I31187,g33498,I31191,I31192,g33499,I31196,I31197,g33500,I31201,I31202,g33501,I31206,
    I31207,g33502,I31211,I31212,g33503,I31216,I31217,g33504,I31221,I31222,g33505,I31226,
    I31227,g33506,I31231,I31232,g33507,I31236,I31237,g33508,I31241,I31242,g33509,I31246,
    I31247,g33510,I31251,I31252,g33511,I31256,I31257,g33512,I31261,I31262,g33513,I31266,
    I31267,g33514,I31271,I31272,g33515,I31276,I31277,g33516,I31281,I31282,g33517,I31286,
    I31287,g33518,I31291,I31292,g33519,I31296,I31297,g33520,I31301,I31302,g33521,I31306,
    I31307,g33522,I31311,I31312,g33523,I31316,I31317,g33524,I31321,I31322,g33525,I31326,
    I31327,g33526,I31331,I31332,g33527,I31336,I31337,g33528,I31341,I31342,g33529,I31346,
    I31347,g33530,I31351,I31352,g33531,I31356,I31357,g33532,g33639,g33640,g33646,g33647,
    g33652,g33657,g33674,g33675,g33676,g33677,g33678,g33680,g33681,g33683,g33684,g33687,
    g33689,g33690,g33693,g33697,g33700,g33701,g33704,g33707,g33710,g33711,g33715,g33717,
    g33718,g33719,g33720,g33721,g33722,g33723,g33724,g33725,g33727,g33728,g33730,g33731,
    I31593,g33734,g33735,I31600,g33742,g33743,g33758,g33759,g33760,g33784,g33785,g33786,
    g33787,g33789,g33790,g33795,g33796,g33798,g33801,g33802,g33803,g33805,g33807,g33808,
    g33809,g33810,g33811,g33812,g33814,g33815,g33816,g33817,g33818,g33819,g33820,g33821,
    g33822,g33828,g33829,g33830,g33831,g33832,g33833,g33834,g33835,g33836,g33837,g33840,
    g33841,g33842,g33843,g33844,g33846,g33847,g33848,g33849,g33855,g33856,g33857,g33858,
    g33859,g33860,g33861,g33862,g33863,g33864,g33865,g33866,g33867,g33868,g33869,g33870,
    g33871,g33872,g33873,g33876,g33877,g33878,g33879,g33880,g33881,g33882,g33883,g33884,
    g33885,g33886,g33887,g33889,g33890,g33892,g33893,g33896,g33897,g33898,g33899,g33900,
    g33901,g33902,g33903,g33904,g33905,g33906,g33907,g33908,g33909,g33910,g33911,g33913,
    g33915,g33919,g33921,g33922,g33924,g33927,g33941,g33942,g33943,g34045,g34050,g34054,
    g34061,g34063,g34065,g34066,g34069,g34071,g34072,g34073,g34074,g34075,g34076,g34077,
    g34078,g34079,g34080,g34081,g34082,g34083,g34084,g34085,g34086,g34087,g34088,g34089,
    g34091,g34092,g34093,g34096,g34097,g34098,g34102,g34104,g34105,g34106,g34108,g34109,
    g34110,g34111,g34112,g34113,g34114,g34115,g34116,g34117,g34119,g34120,g34133,g34135,
    g34136,g34137,g34138,g34139,g34140,g34141,g34143,g34146,g34157,g34169,g34171,g34173,
    g34178,g34179,g34180,g34182,g34183,g34184,g34185,g34186,g34187,g34191,g34196,g34198,
    g34203,g34205,g34211,g34212,g34213,g34214,g34215,g34216,g34217,g34218,g34219,g34223,
    g34224,g34225,g34226,g34228,g34230,g34279,g34281,g34284,g34287,g34291,g34295,g34298,
    g34301,g34309,g34310,g34319,g34322,g34324,g34329,g34333,g34334,g34335,g34337,g34338,
    g34340,g34341,g34342,g34344,g34348,g34363,g34364,g34365,g34367,g34370,g34371,g34375,
    g34378,g34380,g34381,g34382,g34385,g34386,g34388,g34389,g34390,g34393,g34394,g34395,
    g34396,g34397,g34398,g34401,g34410,g34413,g34414,g34415,g34470,g34474,g34475,g34476,
    g34477,g34478,g34479,g34481,g34482,g34483,g34484,g34485,g34486,g34487,g34488,g34489,
    g34492,g34493,g34495,g34497,g34498,g34499,g34500,g34502,g34503,g34506,g34507,g34508,
    g34509,g34513,g34514,g34515,g34516,g34517,g34518,g34519,g34520,g34523,g34524,g34525,
    g34526,g34527,g34528,g34529,g34532,g34533,g34534,g34538,g34541,g34542,g34554,g34555,
    g34556,g34557,g34558,g34560,g34561,g34562,g34563,g34564,g34565,g34566,g34567,g34568,
    g34571,g34572,g34577,g34578,g34580,g34581,g34582,g34584,g34585,g34586,g34588,g34655,
    g34658,g34661,g34662,g34665,g34666,g34667,g34678,g34679,g34681,g34684,g34685,g34686,
    g34687,g34694,g34696,g34700,g34701,g34702,g34706,g34707,g34709,g34710,g34715,g34738,
    g34740,g34741,g34742,g34743,g34744,g34745,g34746,g34747,g34748,g34750,g34751,g34752,
    g34753,g34754,g34756,g34757,g34758,g34763,g34764,g34765,g34771,g34774,g34782,g34811,
    g34841,g34842,g34857,g34858,g34859,g34860,g34861,g34862,g34863,g34865,g34866,g34867,
    g34868,g34869,g34870,g34871,g34872,g34873,g34874,g34875,g34876,g34909,g34948,g34953,
    g34955,g34961,g34962,g34963,g34964,g34965,g34966,g34967,g34968,g34969,g34999,g7404,
    g7450,g7673,g7684,g7764,g7834,g7932,I12583,g8417,g8461,I12611,g8476,g8679,I12782,
    I12783,g8790,g8863,g8904,g8905,I12902,I12903,g8921,g8956,g8957,g9012,g9013,g9055,g9483,
    g9535,g9536,g9984,g10589,g10800,g10802,g11025,g11370,g11372,g11380,g11737,g12768,
    g12911,g12925,g12954,g12981,g12982,g13006,g13077,g13091,g13095,g13155,g13211,g13242,
    g13289,g13295,g13296,g13300,g13385,g13526,g13540,g13543,g13570,g13597,g13623,g13657,
    g13660,g13662,g13699,g13728,g13761,g13762,g13794,g13820,g13858,g13888,g13914,g13938,
    g13941,g13969,g13972,g13973,g13997,g14030,g14044,g14062,g14078,g14119,g14182,g14187,
    g14309,g14387,g14511,g14583,g14844,g14888,g14936,g14977,g15017,g15124,g15125,g15582,
    g15727,g15732,g15789,g15792,g15800,g15803,g15910,g15935,g15965,g15968,g16021,g16022,
    g16052,g16076,g16173,g16187,g16239,g16258,g16261,g16430,g16448,g16506,g16800,g16810,
    g16811,g16839,g16866,g16867,g16876,g16882,g16883,g16926,g16927,g16928,g16959,g16970,
    g17264,g17268,I18385,g17464,I18417,g17488,I18421,g17490,I18449,g17510,I18452,g17511,
    I18492,g17569,I18495,g17570,I18543,g17594,g18879,g18994,g19267,g19274,g19336,g19337,
    g19344,g19356,g19359,g19363,g19441,g19449,g19467,g19475,g19486,g19488,g19501,g19522,
    g19525,g19534,g19535,g19555,g19557,g19572,g19575,g19576,g19587,g19593,g19595,g19604,
    g19605,g19619,g19879,g19904,g19949,g20034,g20051,g20063,g20077,g20082,g20083,g20148,
    g20160,g20169,g20187,g20196,g20202,g20217,g20241,g20276,g20522,g20905,g21891,g21892,
    g21893,g21894,g21895,g21896,g21897,g21898,g21899,g21900,g21901,g22152,g22217,g22225,
    g22226,g22304,g22318,g22331,g22447,g22487,g22490,g22516,g22530,g22531,g22547,g22585,
    g22591,g22625,g22634,g22636,g22639,g22640,g22641,g22644,g22645,g22648,g22652,g22653,
    g22659,g22662,g22664,g22669,g22679,g22684,g22707,g22708,g22751,g22832,g22872,g22901,
    g23087,g23129,g23153,I22267,g23162,g23171,g23183,I22280,g23184,g23193,g23194,g23197,
    I22298,g23198,g23209,g23217,g23251,g23255,g23261,g23262,g23275,g23276,g23296,g23297,
    g23298,g23317,g23318,g23319,g23345,g23346,g23358,g23374,g23383,g23405,g23574,g23615,
    I22830,g23687,g23716,g23720,I22852,g23721,g23750,I22880,g23751,g23770,I22912,g23771,
    g23795,I22958,g23796,g23822,g23825,g23989,g23997,I23162,I23163,g24200,g24201,g24202,
    g24203,g24204,g24205,g24206,g24207,g24208,g24209,g24210,g24211,g24212,g24213,g24214,
    g24215,g24216,g24231,g24232,g24233,g24234,g24235,g24236,g24237,g24238,g24239,g24240,
    g24241,g24242,g24243,g24244,g24245,g24246,g24247,g24248,g24249,g24250,g24251,g24252,
    g24253,g24254,g24255,g24256,g24257,g24258,g24259,g24260,g24261,g24262,g24263,g24264,
    g24265,g24266,g24267,g24268,g24269,g24270,g24271,g24272,g24273,g24274,g24275,g24276,
    g24277,g24278,g24279,g24280,g24281,g24282,g24334,g24335,g24336,g24337,g24338,g24339,
    g24340,g24341,g24342,g24343,g24344,g24345,g24346,g24347,g24348,g24349,g24350,g24351,
    g24352,g24353,g24354,g24355,g24363,g24374,g24390,g24398,g24401,g24430,g24432,g24433,
    g24443,g24444,g24447,g24457,g24460,g24468,g24471,g24478,g24496,g24500,g24510,g24517,
    g24518,g24557,I23755,I23756,g24561,g24565,g24577,g24578,g24580,g24641,g24653,g24705,
    g24715,g24746,g24782,g24799,g24813,g24821,g24840,g24841,g24842,g24853,g24854,g24879,
    g24896,g24907,g24919,g24935,g24946,I24117,g24952,g24965,g24968,g25010,g25037,g25261,
    g25539,g25545,g25575,g25576,g25577,g25591,g25592,g25593,g25594,g25595,g25596,g25597,
    g25598,g25599,g25600,g25601,g25602,g25603,g25604,g25605,g25606,g25607,g25608,g25609,
    g25610,g25611,g25612,g25613,g25614,g25615,g25616,g25617,g25618,g25619,g25621,g25622,
    g25623,g25624,g25625,g25626,g25627,g25628,g25629,g25630,g25631,g25632,g25633,g25634,
    g25635,g25636,g25637,g25638,g25639,g25643,g25644,g25645,g25646,g25647,g25648,g25649,
    g25650,g25651,g25652,g25653,g25654,g25655,g25656,g25657,g25658,g25659,g25660,g25661,
    g25662,g25663,g25664,g25665,g25666,g25667,g25668,g25669,g25670,g25671,g25672,g25673,
    g25674,g25675,g25676,g25677,g25678,g25679,g25680,g25681,g25682,g25683,g25684,g25685,
    g25686,g25687,g25688,g25689,g25690,g25691,g25693,g25694,g25695,g25696,g25697,g25698,
    g25699,g25700,g25701,g25702,g25703,g25704,g25705,g25706,g25707,g25708,g25709,g25710,
    g25711,g25712,g25713,g25714,g25715,g25716,g25717,g25718,g25719,g25720,g25721,g25722,
    g25723,g25724,g25725,g25726,g25727,g25728,g25729,g25730,g25731,g25732,g25733,g25734,
    g25735,g25736,g25737,g25738,g25739,g25740,g25741,g25742,g25743,g25744,g25745,g25746,
    g25747,g25748,g25749,g25750,g25751,g25752,g25753,g25754,g25755,g25756,g25757,g25758,
    g25759,g25760,g25761,g25762,g25763,g25764,g25767,g25774,g25789,g25791,g25805,g25819,
    g25821,g25834,g25835,g25836,g25839,g25856,g25867,g25868,g25877,g25878,g25885,g25894,
    g25906,g25910,g25911,g25917,g25929,g25935,g25936,g25937,g25940,g25941,g25942,g25943,
    g25945,g25960,g26080,g26082,g26089,g26099,g26278,g26293,g26299,g26305,g26327,g26328,
    g26329,g26334,g26335,g26342,g26343,g26344,g26348,g26349,g26359,g26361,g26363,g26365,
    g26377,g26386,g26392,g26396,g26422,g26512,g26616,g26636,g26657,g26673,g26690,g26694,
    g26703,g26721,g26725,g26733,g26737,g26751,g26755,g26759,g26766,g26770,g26781,g26785,
    g26789,g26793,g26800,g26805,g26809,g26813,g26866,I25612,I25613,g26874,g26878,g26879,
    g26880,g26881,g26882,g26883,g26884,g26885,g26886,g26887,g26888,g26889,g26890,g26891,
    g26892,g26893,g26894,g26895,g26896,g26897,g26898,g26899,g26900,g26901,g26902,g26903,
    g26904,g26905,g26906,g26907,g26908,g26909,g26910,g26911,g26912,g26913,g26914,g26915,
    g26916,g26917,g26918,g26919,g26920,g26921,g26922,g26923,g26924,g26925,g26926,g26927,
    g26928,g26929,g26930,g26931,g26932,g26933,g26934,g26938,g26939,g26940,g26944,g26945,
    g26946,g26947,g26948,g26949,g26950,g26951,g26952,g26953,g26954,g26955,g26956,g26957,
    g26958,g26959,g26960,g26961,g26962,g26963,g26964,g26965,g26966,g26967,g26968,g26969,
    g26970,g26971,g26972,I25736,g27008,g27016,g27019,g27024,g27026,g27031,g27037,g27108,
    g27122,g27126,g27133,g27135,g27147,g27150,g27152,g27159,g27179,g27182,g27205,g27224,
    g27225,g27226,g27231,g27232,g27233,g27236,g27238,g27239,g27240,g27241,g27243,g27244,
    g27248,g27250,g27253,g27257,g27258,g27261,g27271,g27274,g27278,g27283,g27289,g27290,
    g27383,g27394,g27403,g27405,g27426,g27429,g27431,g27450,g27453,g27456,g27458,g27484,
    g27487,g27489,g27506,g27509,g27515,g27524,g27532,g27533,g27542,g27543,g27544,g27551,
    g27552,g27555,g27556,g27561,g27562,g27563,g27566,g27567,g27569,g27570,g27571,g27572,
    g27574,g27575,g27578,g27579,g27580,g27581,g27584,g27589,g27590,g27591,g27596,g27663,
    g27742,g27779,g27800,g27837,g27858,g27886,g27907,g27937,g27970,g27972,g27974,g27980,
    I26522,I26523,g28043,g28044,g28045,g28046,g28047,g28048,g28049,g28050,g28051,g28052,
    g28053,g28054,g28055,g28056,g28057,g28058,g28059,g28060,g28061,g28062,g28063,g28064,
    g28065,g28066,g28067,g28068,g28069,g28070,g28071,g28072,g28073,g28074,g28075,g28076,
    g28077,g28078,g28082,g28083,g28084,g28085,g28086,g28087,g28088,g28089,g28090,g28091,
    g28092,g28093,g28094,g28095,g28096,g28097,g28098,g28099,g28100,g28101,g28102,g28103,
    g28104,g28105,g28118,g28132,g28134,g28135,g28138,I26643,I26644,g28140,g28172,g28179,
    g28180,g28186,g28188,g28191,g28194,g28208,g28209,g28211,g28212,g28216,I26741,I26742,
    g28220,g28230,g28279,g28286,g28295,g28296,g28297,g28305,g28306,g28308,g28309,g28310,
    g28316,g28317,g28319,g28320,g28322,g28323,g28328,g28329,g28331,g28332,g28334,g28335,
    g28342,g28344,g28345,g28347,g28348,g28357,g28358,g28359,g28361,g28362,g28368,g28369,
    g28371,g28372,g28373,g28374,g28375,g28385,g28386,g28387,g28388,g28389,g28390,g28400,
    g28401,g28402,g28403,g28404,g28405,g28416,g28417,g28418,g28419,g28420,g28428,g28429,
    g28430,g28435,g28490,g28497,g28511,g28513,g28517,g28518,g28525,g28526,g28527,g28533,
    g28534,g28536,g28538,g28544,g28545,g28546,g28548,g28549,g28551,g28560,g28561,g28562,
    g28564,g28565,g28566,g28574,g28576,g28577,g28578,g28580,g28581,g28582,g28589,g28591,
    g28592,g28594,g28595,g28596,g28600,g28603,g28605,g28607,g28609,g28610,g28611,g28613,
    g28614,g28618,g28619,g28621,g28622,g28623,g28625,g28628,g28629,g28631,g28632,g28634,
    g28635,g28636,g28640,g28641,g28643,g28644,g28646,g28647,g28649,g28650,g28651,g28659,
    g28661,g28662,g28664,g28665,g28667,g28668,g28670,g28671,g28680,g28681,g28682,g28684,
    g28685,g28687,g28688,g28690,g28691,g28698,g28699,g28700,g28701,g28702,g28704,g28705,
    g28707,g28708,g28715,g28716,g28717,g28718,g28719,g28720,g28721,g28723,g28724,g28727,
    g28728,g28729,g28730,g28731,g28732,g28733,g28734,g28735,g28743,g28744,g28745,g28746,
    g28747,g28748,g28749,g28750,g28751,g28772,g28773,g28774,g28775,g28776,g28777,g28778,
    g28814,g28815,g28816,g28817,g28818,g28850,g28851,g28852,g28884,g29068,g29078,g29105,
    g29114,g29143,g29148,g29166,g29168,g29176,g29197,g29222,g29223,g29224,g29225,g29226,
    g29227,g29228,g29229,g29230,g29231,g29232,g29233,g29234,g29235,g29236,g29237,g29238,
    g29239,g29240,g29241,g29242,g29243,g29244,g29245,g29246,g29247,g29248,g29249,g29250,
    g29251,g29252,g29253,g29254,g29255,g29256,g29257,g29258,g29259,g29260,g29261,g29262,
    g29263,g29264,g29265,g29266,g29267,g29268,g29269,g29270,g29271,g29272,g29273,g29274,
    g29275,g29276,g29277,g29278,g29279,g29280,g29281,g29282,g29283,g29284,g29285,g29286,
    g29287,g29288,g29289,g29290,g29291,g29292,g29293,g29294,g29295,g29296,g29297,g29298,
    g29299,g29300,g29301,g29302,g29303,g29304,g29305,g29306,g29307,g29308,g29309,g29313,
    g29319,g29325,g29366,g29373,g29476,g29478,g29479,g29480,g29481,g29482,g29483,g29484,
    g29485,g29486,g29487,g29488,g29489,g29490,g29495,g29496,g29501,g29502,g29504,g29506,
    g29508,g29520,g29529,g29539,g29583,g29643,g29692,g29706,g29716,g29717,g29730,g29734,
    g29735,g29741,g29748,g29753,g29754,g29756,g29763,g29764,g29768,g29775,g29776,g29777,
    g29786,g29790,g29791,g29792,g29793,g29801,g29802,g29813,g29848,g29849,g29864,g29879,
    g29892,g29904,I28147,g29914,g30081,g30092,g30093,g30103,g30104,g30114,g30115,g30127,
    g30128,g30141,g30163,g30176,g30189,g30201,g30214,g30270,g30279,g30286,g30287,g30291,
    g30293,g30298,g30300,g30304,g30307,g30311,g30314,I28566,I28567,g30317,g30333,g30334,
    g30335,g30336,g30337,g30338,g30339,g30340,g30341,g30342,g30343,g30344,g30345,g30346,
    g30347,g30348,g30349,g30350,g30351,g30352,g30353,g30354,g30355,g30356,g30357,g30358,
    g30359,g30360,g30361,g30362,g30363,g30364,g30365,g30366,g30367,g30368,g30369,g30370,
    g30371,g30372,g30373,g30374,g30375,g30376,g30377,g30378,g30379,g30380,g30381,g30382,
    g30383,g30384,g30385,g30386,g30387,g30388,g30389,g30390,g30391,g30392,g30393,g30394,
    g30395,g30396,g30397,g30398,g30399,g30400,g30401,g30402,g30403,g30404,g30405,g30406,
    g30407,g30408,g30409,g30410,g30411,g30412,g30413,g30414,g30415,g30416,g30417,g30418,
    g30419,g30420,g30421,g30422,g30423,g30424,g30425,g30426,g30427,g30428,g30429,g30430,
    g30431,g30432,g30433,g30434,g30435,g30436,g30437,g30438,g30439,g30440,g30441,g30442,
    g30443,g30444,g30445,g30446,g30447,g30448,g30449,g30450,g30451,g30452,g30453,g30454,
    g30455,g30456,g30457,g30458,g30459,g30460,g30461,g30462,g30463,g30464,g30465,g30466,
    g30467,g30468,g30469,g30470,g30471,g30472,g30473,g30474,g30475,g30476,g30477,g30478,
    g30479,g30480,g30481,g30482,g30483,g30484,g30485,g30486,g30487,g30488,g30489,g30490,
    g30491,g30492,g30493,g30494,g30495,g30496,g30497,g30498,g30499,g30500,g30501,g30502,
    g30503,g30504,g30505,g30506,g30507,g30508,g30509,g30510,g30511,g30512,g30513,g30514,
    g30515,g30516,g30517,g30518,g30519,g30520,g30521,g30522,g30523,g30524,g30525,g30526,
    g30527,g30528,g30529,g30530,g30531,g30532,g30533,g30534,g30535,g30536,g30537,g30538,
    g30539,g30540,g30541,g30542,g30543,g30544,g30545,g30546,g30547,g30548,g30549,g30550,
    g30551,g30552,g30553,g30554,g30555,g30556,g30557,g30558,g30559,g30560,g30561,g30562,
    g30563,g30579,g30597,g30605,g30608,g30609,g30611,g30672,g30732,g30733,g30734,g30824,
    g30916,g30984,g31001,g31002,g31007,g31014,g31020,g31144,g31221,g31241,g31244,g31245,
    g31246,g31247,g31248,g31249,g31250,g31251,g31253,g31254,g31255,g31256,g31257,g31258,
    g31259,g31260,g31267,g31268,g31269,g31274,g31276,g31277,g31279,g31284,g31287,g31288,
    g31289,g31291,g31293,g31295,g31302,g31303,g31304,g31306,g31307,g31308,g31311,g31315,
    g31316,g31317,g31319,g31320,g31322,g31325,g31326,g31375,g31465,g31466,g31468,g31472,
    g31473,g31474,g31591,g31668,g31670,g31745,g31749,g31751,g31754,g31755,g31757,g31760,
    g31761,g31762,g31764,g31766,g31767,g31768,g31770,g31772,g31773,g31774,g31775,g31779,
    g31781,g31782,I29351,I29352,g31783,g31785,g31864,g31865,g31866,g31867,g31868,g31869,
    g31870,g31871,g31872,g31873,g31874,g31875,g31876,g31877,g31878,g31879,g31880,g31881,
    g31882,g31883,g31884,g31885,g31886,g31887,g31888,g31889,g31890,g31891,g31892,g31893,
    g31894,g31895,g31896,g31897,g31898,g31899,g31900,g31901,g31902,g31903,g31904,g31905,
    g31906,g31907,g31908,g31909,g31910,g31911,g31912,g31913,g31914,g31915,g31916,g31917,
    g31918,g31919,g31920,g31921,g31922,g31923,g31924,g31925,g31926,g31927,g31928,g31929,
    g31930,g31931,g31932,g31964,g32037,g32094,g32117,g32123,g32124,g32125,g32130,g32131,
    g32132,g32144,g32155,g32202,g32208,g32209,g32210,g32211,g32216,g32217,g32218,g32219,
    g32220,g32221,g32222,g32223,g32225,g32226,g32227,g32228,g32229,g32230,g32231,g32233,
    g32235,g32236,g32237,g32238,g32239,g32240,g32243,g32245,g32247,g32249,g32250,g32251,
    g32252,g32253,g32257,g32259,g32262,g32264,g32266,g32267,g32268,g32271,g32275,g32277,
    g32279,g32280,g32285,g32288,g32289,g32294,g32344,g32346,g32347,g32349,g32351,g32352,
    g32353,g32354,g32355,g32357,g32358,g32359,g32360,g32361,g32362,g32367,g32368,g32370,
    g32371,g32372,g32373,g32374,g32375,g32380,g32385,g32386,g32387,g32388,g32389,g32390,
    g32391,g32392,g32395,g32398,g32399,g32408,g32426,g32427,I29985,I29986,I30054,I30055,
    I30123,I30124,I30192,I30193,I30261,I30262,I30330,I30331,I30399,I30400,I30468,I30469,
    g32976,g32977,g32978,g32979,g32980,g32981,g32982,g32983,g32984,g32985,g32986,g32987,
    g32988,g32989,g32990,g32991,g32992,g32993,g32994,g32995,g32996,g32997,g32998,g32999,
    g33000,g33001,g33002,g33003,g33004,g33005,g33006,g33007,g33008,g33009,g33010,g33011,
    g33012,g33013,g33014,g33015,g33016,g33017,g33018,g33019,g33020,g33021,g33022,g33023,
    g33024,g33025,g33026,g33027,g33028,g33029,g33030,g33031,g33032,g33033,g33034,g33035,
    g33036,g33037,g33038,g33039,g33040,g33041,g33042,g33043,g33044,g33045,g33046,g33047,
    g33048,g33049,g33050,g33051,g33052,g33053,g33054,g33055,g33056,g33057,g33058,g33059,
    g33060,g33061,g33062,g33063,g33064,g33065,g33066,g33067,g33068,g33069,g33070,g33076,
    g33115,g33116,g33118,g33119,g33123,I30717,I30718,g33149,g33159,I30727,I30728,g33164,
    I30734,I30735,g33176,I30740,I30741,g33187,I30745,I30746,g33197,I30750,I30751,g33204,
    I30755,I30756,g33212,I30760,I30761,g33219,g33227,g33231,g33232,g33234,g33235,g33236,
    g33238,g33240,g33251,g33253,g33254,g33255,g33256,g33257,g33259,g33260,g33261,g33262,
    g33265,g33266,g33267,g33268,g33270,g33271,g33272,g33273,g33274,g33275,g33276,g33277,
    g33278,g33279,g33280,g33281,g33282,g33283,g33286,g33287,g33288,g33289,g33290,g33291,
    g33292,g33293,g33294,g33295,g33296,g33297,g33298,g33303,g33310,g33312,g33313,g33314,
    g33315,g33316,g33317,g33318,g33321,g33323,g33380,g33383,g33384,g33386,g33387,g33389,
    g33390,g33393,g33534,g33535,g33536,g33537,g33538,g33539,g33540,g33541,g33542,g33543,
    g33544,g33545,g33546,g33547,g33548,g33549,g33550,g33551,g33552,g33553,g33554,g33555,
    g33556,g33557,g33558,g33559,g33560,g33561,g33562,g33563,g33564,g33565,g33566,g33567,
    g33568,g33569,g33570,g33571,g33572,g33573,g33574,g33575,g33576,g33577,g33578,g33579,
    g33580,g33581,g33582,g33583,g33584,g33585,g33586,g33587,g33588,g33589,g33590,g33591,
    g33592,g33593,g33594,g33595,g33596,g33597,g33598,g33599,g33600,g33601,g33602,g33603,
    g33604,g33605,g33606,g33607,g33608,g33609,g33610,g33611,g33612,g33613,g33614,g33615,
    g33616,g33617,g33618,g33619,g33620,g33621,g33622,g33623,g33624,g33625,g33626,g33627,
    g33628,g33685,g33692,g33694,g33699,g33703,g33706,g33709,g33714,g33732,g33733,g33788,
    g33791,g33794,g33891,g33914,I31838,I31839,g33951,I31843,I31844,g33952,I31848,I31849,
    g33953,I31853,I31854,g33954,I31858,I31859,g33955,I31863,I31864,g33956,I31868,I31869,
    g33957,I31873,I31874,g33958,g33960,g33961,g33962,g33963,g33964,g33965,g33966,g33967,
    g33968,g33969,g33970,g33971,g33972,g33973,g33974,g33975,g33976,g33977,g33978,g33979,
    g33980,g33981,g33982,g33983,g33984,g33985,g33986,g33987,g33988,g33989,g33990,g33991,
    g33992,g33993,g33994,g33995,g33996,g33997,g33998,g33999,g34000,g34001,g34002,g34003,
    g34004,g34005,g34006,g34007,g34008,g34009,g34010,g34011,g34012,g34013,g34014,g34015,
    g34016,g34017,g34018,g34019,g34020,g34021,g34022,g34023,g34024,g34025,g34026,g34027,
    g34028,g34029,g34030,g34031,g34032,g34033,g34034,g34035,g34036,g34037,g34038,g34039,
    g34040,g34041,g34043,g34046,g34055,g34057,g34064,g34090,g34095,g34099,g34100,g34101,
    g34103,g34107,g34125,g34127,g34148,g34149,g34153,g34158,g34166,g34167,g34168,g34170,
    g34172,g34189,g34190,g34193,g34194,g34199,g34204,g34206,g34207,g34231,g34249,g34250,
    g34251,g34252,g34253,g34254,g34255,g34256,g34257,g34258,g34259,g34260,g34261,g34262,
    g34263,g34264,g34265,g34266,g34267,g34268,g34269,g34273,g34274,g34278,g34280,g34282,
    g34283,g34286,g34288,g34289,g34290,g34292,g34293,g34294,g34297,g34300,g34303,g34305,
    g34306,g34314,g34318,g34321,g34330,g34331,g34332,g34347,g34349,g34350,g34352,g34353,
    g34366,g34368,g34369,g34372,g34373,g34374,g34376,g34377,g34379,g34399,g34402,g34403,
    g34404,g34405,g34406,g34407,g34411,g34412,g34416,g34417,g34421,g34438,g34439,g34440,
    g34441,g34442,g34443,g34444,g34445,g34446,g34447,g34448,g34449,g34450,g34451,g34452,
    g34453,g34454,g34455,g34456,g34457,g34458,g34459,g34460,g34461,g34462,g34463,g34464,
    g34465,g34466,g34467,g34468,g34494,g34535,g34537,g34598,g34599,g34600,g34601,g34602,
    g34603,g34604,g34605,g34606,g34607,g34608,g34609,g34610,g34611,g34612,g34613,g34614,
    g34615,g34616,g34617,g34618,g34619,g34620,g34621,g34622,g34623,g34624,g34625,g34626,
    g34627,g34628,g34629,g34630,g34631,g34632,g34633,g34634,g34635,g34636,g34637,g34638,
    g34639,g34640,g34641,g34642,g34643,g34644,g34645,g34646,g34647,g34649,g34657,g34663,
    g34693,g34695,g34708,g34719,g34720,g34721,g34722,g34723,g34724,g34725,g34726,g34727,
    g34728,g34729,g34730,g34731,g34732,g34733,g34734,g34735,g34761,g34762,g34781,g34783,
    g34790,g34791,g34792,g34793,g34794,g34795,g34796,g34797,g34798,g34799,g34800,g34801,
    g34802,g34803,g34804,g34805,g34806,g34807,g34808,g34809,g34819,g34826,g34843,g34849,
    g34850,g34856,g34880,g34881,g34882,g34884,g34887,g34890,g34894,g34897,g34900,g34903,
    g34906,g34911,g34931,g34957,g34970,g34971,g34974,g34975,g34976,g34977,g34978,g34979,
    g34980,g35000,I11824,I11825,I11826,g7133,g7150,g7167,g7184,I11864,I11865,I11866,g7201,
    g7209,I11877,I11878,I11879,g7223,g7227,g7228,g7442,g7549,g7582,I12074,I12075,I12076,
    g7598,g7611,I12096,I12097,I12098,g7620,g7690,g7701,I12203,I12204,I12205,g7803,I12217,
    I12218,I12219,g7823,g7836,g7846,g7850,I12240,I12241,I12242,g7857,I12251,I12252,I12253,
    g7869,I12261,I12262,I12263,g7879,I12269,I12270,I12271,g7885,I12277,I12278,I12279,
    g7887,I12287,I12288,I12289,g7897,I12344,I12345,I12346,g8010,I12372,I12373,I12374,
    g8069,g8105,I12401,I12402,I12403,g8124,g8163,g8227,I12468,I12469,I12470,g8238,g8292,
    g8347,I12544,I12545,I12546,g8359,g8434,g8500,g8561,g8609,g8632,g8678,g8691,g8728,
    I12728,I12729,I12730,g8737,g8751,g8769,g8803,g8806,g8829,g8847,I12840,I12841,I12842,
    g8871,I12848,I12849,I12850,g8873,g8889,I12876,I12877,I12878,g8913,g8967,g9092,g9177,
    g9203,g9246,I13043,I13044,I13045,g9258,I13065,I13066,I13067,g9295,I13077,I13078,
    I13079,g9310,g9334,g9372,I13109,I13110,I13111,g9391,g9442,I13139,I13140,I13141,g9461,
    g9485,g9509,I13182,I13183,I13184,g9528,g9538,g9543,g9567,g9591,g9595,g9629,g9645,g9654,
    g9663,g9705,g9715,g9724,I13334,I13335,I13336,g9750,g9775,g9800,I13382,I13383,I13384,
    g9823,I13390,I13391,I13392,g9825,I13401,I13402,I13403,g9830,g9852,g9883,I13442,I13443,
    I13444,g9904,I13452,I13453,I13454,g9908,I13462,I13463,I13464,g9912,g9954,I13497,I13498,
    I13499,g9966,I13509,I13510,I13511,g9972,I13518,I13519,I13520,g9975,g10022,I13564,
    I13565,I13566,g10041,g10124,g10160,g10185,g10207,g10224,I13729,I13730,I13731,g10307,
    I13749,I13750,I13751,g10336,I13850,I13851,I13852,g10472,g10511,g10515,g10520,g10529,
    g10537,g10550,g10551,g10552,g10556,g10561,g10566,g10567,g10568,g10569,g10573,g10578,
    g10583,g10584,g10585,g10586,g10587,g10598,g10601,g10602,g10603,g10604,g10605,g10609,
    g10610,g10611,g10614,g10617,g10618,g10622,g10623,g10653,g10726,g10737,g10738,g10754,
    g10755,g10759,g10775,g10796,g10820,g10905,g10909,g10916,g10928,g10929,g10935,g10939,
    g10946,g10951,g10961,g10971,g11002,g11020,g11117,I14169,I14170,I14171,g11118,g11130,
    g11134,I14185,I14186,I14187,g11135,g11149,I14204,I14205,I14206,g11153,I14211,I14212,
    I14213,g11154,g11155,I14228,I14229,I14230,g11169,g11172,g11173,I14247,I14248,I14249,
    g11189,g11190,I14257,I14258,I14259,g11193,g11200,I14275,I14276,I14277,g11206,I14289,
    I14290,I14291,g11224,g11245,g11251,g11279,I14330,I14331,I14332,g11292,g11302,g11312,
    g11320,I14350,I14351,I14352,g11323,g11326,g11330,I14368,I14369,I14370,g11350,g11355,
    g11356,g11374,g11381,g11382,I14398,I14399,I14400,g11389,g11394,g11395,g11396,g11405,
    g11409,g11410,g11411,g11412,I14427,I14428,I14429,g11419,g11424,g11426,g11432,g11441,
    g11442,g11443,g11444,g11445,g11446,g11479,g11480,g11489,g11490,g11491,g11492,I14480,
    I14481,I14482,g11511,g11533,g11534,g11543,g11544,I14497,I14498,I14499,g11545,I14508,
    I14509,I14510,g11559,I14516,I14517,I14518,g11561,g11590,I14530,I14531,I14532,g11591,
    g11639,g11674,g11675,g11676,g11679,g11707,g11708,I14609,I14610,I14611,g11761,g11858,
    g11881,g11892,g11903,I14712,I14713,I14714,g11906,g11914,I14733,I14734,I14735,g11923,
    g11933,g11934,g11936,g11938,I14764,I14765,I14766,g11944,g11951,g11952,g11953,g11955,
    g11957,g11959,g11961,I14788,I14789,I14790,g11962,g11968,g11969,g11970,g11971,g11973,
    g11974,g11975,g11977,g11979,I14816,I14817,I14818,g11980,g11990,g11992,g11993,g11994,
    g11996,g11997,g11998,g12000,I14853,I14854,I14855,g12001,g12008,g12014,g12016,g12019,
    g12020,g12022,g12023,g12024,I14883,I14884,I14885,g12028,g12035,g12042,g12044,g12045,
    g12048,g12049,g12052,g12053,I14923,I14924,I14925,g12066,g12073,g12078,g12079,g12080,
    g12083,g12084,g12087,I14955,I14956,I14957,g12100,g12111,g12112,g12114,g12115,g12116,
    g12118,g12119,g12120,g12124,g12125,I14991,I14992,I14993,g12136,I15002,I15003,I15004,
    g12144,g12145,g12147,g12148,g12149,g12151,g12152,g12153,g12155,g12159,g12169,g12185,
    I15041,I15042,I15043,g12187,g12188,g12190,I15051,I15052,I15053,g12191,g12192,g12194,
    g12195,g12196,g12197,g12207,I15078,I15079,I15080,g12221,g12222,I15087,I15088,I15089,
    g12224,g12225,g12227,g12232,I15105,I15106,I15107,g12239,g12244,g12245,g12255,I15121,
    I15122,I15123,g12285,I15128,I15129,I15130,g12286,g12287,g12289,g12292,g12293,g12294,
    I15147,I15148,I15149,g12301,g12306,g12307,g12317,g12323,I15166,I15167,I15168,g12332,
    I15174,I15175,I15176,g12336,g12340,g12341,g12342,g12343,g12344,I15193,I15194,I15195,
    g12351,g12356,g12357,g12369,I15212,I15213,I15214,g12370,g12402,g12411,g12412,g12413,
    g12414,g12415,g12416,I15241,I15242,I15243,g12423,g12428,g12429,I15253,I15254,I15255,
    g12431,I15262,I15263,I15264,g12436,g12449,g12450,g12459,g12460,g12461,g12462,g12463,
    g12464,I15287,I15288,I15289,g12471,g12476,I15298,I15299,I15300,g12478,I15306,I15307,
    I15308,g12482,g12491,g12511,g12512,g12521,g12522,g12523,g12524,g12525,g12526,I15333,
    I15334,I15335,g12538,I15340,I15341,I15342,g12539,g12577,g12578,g12587,g12588,g12589,
    g12590,I15363,I15364,I15365,g12592,g12628,g12629,g12638,g12639,g12644,g12686,g12767,
    g12796,g12797,g12819,g12822,g12910,g12915,g12933,g12941,g12947,g12969,g12971,g12972,
    g12999,g13000,g13040,g13043,g13050,g13057,g13058,g13066,g13067,g13069,g13079,g13083,
    g13084,g13086,g13092,g13093,g13097,g13098,g13100,g13102,g13104,g13105,g13108,g13109,
    g13115,g13118,g13119,g13121,g13124,g13130,g13131,g13134,g13137,g13139,g13143,g13176,
    g13210,g13217,g13240,g13241,g13248,g13256,g13257,g13260,g13264,g13266,g13273,g13281,
    g13283,g13284,g13288,g13291,g13307,g13315,g13330,g13346,g13432,g13459,g13462,g13464,
    g13469,g13475,g13476,g13478,g13479,g13486,g13495,g13496,g13498,g13499,g13511,g13513,
    g13515,g13516,g13527,g13528,g13529,g13544,g13551,g13554,g13573,g13580,g13600,g13627,
    g13628,g13634,g13666,g13667,g13672,g13676,g13708,g13709,g13712,g13727,g13739,g13742,
    g13756,g13764,g13779,g13795,g13797,g13798,g13821,g13822,g13823,g13834,g13846,g13850,
    g13851,g13854,g13855,g13861,g13866,g13867,g13870,g13871,g13873,g13882,g13884,g13886,
    g13889,g13892,g13896,g13897,g13898,g13907,g13909,g13911,g13915,g13918,g13920,g13923,
    g13927,g13928,g13929,g13940,g13945,g13948,g13951,g13955,g13958,g13960,g13963,g13967,
    g13968,g13977,g13980,g13983,g13986,g13990,g13993,g14005,g14008,g14011,g14014,g14015,
    g14018,g14021,g14024,g14038,g14041,g14045,g14048,g14051,g14054,g14055,g14058,g14066,
    g14069,g14072,g14075,g14079,g14082,g14085,g14088,g14089,g14098,g14101,g14104,g14107,
    g14110,g14113,g14116,g14120,g14123,g14127,g14130,g14133,g14136,g14139,g14142,g14146,
    g14151,g14154,g14157,g14160,g14170,g14177,g14223,g14234,g14254,g14258,g14279,g14317,
    g14333,g14343,g14344,g14378,g14379,g14407,g14408,g14422,g14433,g14434,g14452,g14489,
    g14505,g14517,g14519,g14520,g14521,g14542,g14546,g14547,g14548,g14569,g14570,g14572,
    g14573,g14574,g14590,g14596,g14598,g14599,g14600,g14601,g14625,g14626,g14627,g14636,
    g14637,g14638,g14655,g14656,g14659,g14663,g14664,g14665,g14674,g14675,I16778,I16779,
    I16780,g14677,g14682,g14683,g14686,g14688,g14691,g14695,g14696,g14697,g14706,g14720,
    g14723,g14727,g14730,g14732,g14735,g14739,g14740,g14741,g14750,g14755,g14758,g14761,
    g14764,g14768,g14771,g14773,g14776,g14780,g14781,g14782,g14794,g14797,g14800,g14803,
    g14804,g14807,g14810,g14813,g14817,g14820,g14822,g14825,g14829,g14830,g14838,g14841,
    g14845,g14848,g14851,g14854,g14855,g14858,g14861,g14864,g14868,g14871,g14876,g14879,
    g14882,g14885,g14889,g14892,g14895,g14898,g14899,g14902,g14905,g14908,g14915,g14918,
    g14921,g14924,g14927,g14930,g14933,g14937,g14940,g14943,g14946,g14947,g14950,g14953,
    g14956,g14959,g14962,g14965,g14968,g14971,g14974,g14978,g14981,g14984,g14987,g14993,
    g14996,g14999,g15002,g15005,g15008,g15011,g15014,g15018,g15021,g15024,g15027,g15030,
    g15033,g15036,g15039,g15042,g15045,g15572,g15581,g15591,g15674,g15695,g15702,g15708,
    g15709,g15710,g15713,g15715,g15717,g15719,g15720,g15721,g15723,g15725,g15726,g15728,
    g15729,g15730,g15734,g15735,g15736,g15737,g15741,g15742,g15743,g15744,g15748,g15751,
    g15752,g15753,g15780,g15781,g15782,g15787,g15788,g15798,g15829,g15832,g15833,g15843,
    g15844,g15853,g15864,g15867,g15877,I17379,I17380,I17381,g15904,g15907,I17404,I17405,
    I17406,g15959,g15962,I17446,I17447,I17448,g16069,I17460,I17461,I17462,g16093,g16097,
    I17474,I17475,I17476,g16119,I17494,I17495,I17496,g16155,g16181,g16196,g16225,g16236,
    g16238,g16259,g16260,g16264,g16275,g16278,g16281,g16282,g16291,g16296,g16299,g16304,
    g16306,g16312,g16316,g16319,g16321,g16507,g16524,g16586,g16604,g16625,g16628,g16657,
    g16660,g16663,I17883,I17884,I17885,g16681,g16687,g16694,g16696,I17923,I17924,I17925,
    g16713,g16719,g16723,g16728,g16741,g16745,g16749,g16757,g16770,g16772,g16776,g16813,
    g16815,g16854,g16875,g16893,g16925,g16956,g17137,g17217,g17220,g17225,g17243,g17246,
    g17287,g17290,g17297,g17312,g17315,g17363,g17364,g17396,g17399,g17412,g17468,g17474,
    g17492,g17493,g17495,g17500,g17513,g17514,g17520,g17525,I18485,I18486,I18487,g17568,
    g17571,g17572,g17578,g17581,g17586,I18529,I18530,I18531,g17592,I18536,I18537,I18538,
    g17593,g17595,g17596,g17597,g17598,g17605,g17608,I18579,I18580,I18581,g17618,I18587,
    I18588,I18589,g17624,g17634,g17635,g17640,g17647,g17650,I18625,I18626,I18627,g17656,
    I18633,I18634,I18635,g17662,g17668,g17669,g17670,g17675,g17679,g17686,g17689,I18680,
    I18681,I18682,g17699,g17705,g17706,g17708,g17712,g17716,g17723,g17732,g17734,g17736,
    g17740,g17744,g17748,g17755,g17757,g17761,g17765,g17773,g17775,g17779,g17788,g17790,
    g17792,g17814,g17816,g17820,g17846,g17872,g19265,g19335,g19358,g19442,g19450,g19455,
    g19466,g19474,g19483,g19495,g19506,g19510,g19513,g19530,g19546,g19549,g19589,g19597,
    g19611,g19614,g19632,I20165,I20166,I20167,g19764,I20187,I20188,I20189,g19782,I20203,
    I20204,I20205,g19792,g19795,I20221,I20222,I20223,g19854,g19856,g19857,g19874,g19875,
    g19886,g19903,g19913,g19916,g19962,g19965,g20007,g20011,g20039,g20055,g20068,g20076,
    g20081,g20092,g20107,g20111,g20133,g20134,g20150,g20151,g20161,g20163,g20170,g20172,
    g20173,g20181,g20184,g20185,g20186,g20198,g20199,I20460,I20461,I20462,g20200,I20467,
    I20468,I20469,g20201,g20214,I20486,I20487,I20488,g20216,g20236,g20248,g20271,g20371,
    g20619,g20644,g20645,g20675,g20676,g20733,g20734,g20783,g20784,g20838,g20870,g20871,
    g20979,g21011,g21124,g21186,g21187,g21190,g21253,g21272,g21283,g21287,g21288,g21289,
    g21294,g21301,g21307,g21330,g21331,g21334,g21338,g21339,g21344,g21345,g21350,g21351,
    g21353,g21354,g21356,g21357,g21359,g21360,g21363,g21364,g21365,g21377,g21384,g21385,
    g21386,g21388,g21401,g21402,g21403,g21415,g21416,g21417,g21429,g21432,g21433,g21459,
    g21462,g21509,g21555,g21603,g22306,g22312,g22325,g22638,g22642,g22643,g22650,g22651,
    g22661,I21976,I21977,I21978,g22663,g22666,g22668,I21992,I21993,I21994,g22681,g22687,
    g22688,g22709,g22711,g22712,g22713,g22715,g22753,g22754,g22755,g22757,g22833,g22836,
    g22837,g22838,g22839,g22850,g22852,g22853,g22864,g22874,g22875,g22885,g22902,g22908,
    g22921,g22940,g22941,g22984,g23010,g23047,g23067,g23105,g23112,g23132,g23139,g23167,
    g23195,g23210,g23266,g23281,g23286,g23309,g23324,g23342,g23357,g23379,g23428,I22683,
    I22684,I22685,g23552,I22710,I22711,I22712,g23575,I22717,I22718,I22719,g23576,g23590,
    I22753,I22754,I22755,g23616,I22760,I22761,I22762,g23617,g23623,g23630,I22792,I22793,
    I22794,g23655,I22799,I22800,I22801,g23656,g23659,g23666,I22822,I22823,I22824,g23685,
    g23692,g23699,I22844,I22845,I22846,g23719,g23726,g23733,I22864,I22865,I22866,g23747,
    I22871,I22872,I22873,g23748,g23756,I22892,I22893,I22894,g23761,I22899,I22900,I22901,
    g23762,I22921,I22922,I22923,g23778,I22929,I22930,I22931,g23780,I22936,I22937,I22938,
    g23781,g23782,I22944,I22945,I22946,g23786,I22965,I22966,I22967,g23809,I22972,I22973,
    I22974,g23810,g23850,g23890,g23909,g23932,g23949,g23972,I23118,I23119,I23120,g23975,
    g23978,g24362,I23585,I23586,I23587,g24369,I23600,I23601,I23602,g24380,g24528,g24544,
    g24547,g24566,g24567,g24570,g24574,g24576,g24583,g24584,g24591,g24601,g24609,g24620,
    g24621,g24652,g24661,g24662,g24677,g24678,I23917,I23918,I23919,g24760,g24776,g24787,
    I23949,I23950,I23951,g24792,g24793,I23961,I23962,I23963,g24798,I23969,I23970,I23971,
    g24802,g24804,I23978,I23979,I23980,g24807,I23985,I23986,I23987,g24808,g24809,g24814,
    g24880,g24890,g24905,g24906,g24916,g24917,g24918,g24924,g24925,g24926,g24932,g24933,
    g24934,g24936,g24942,g24943,g24944,g24950,g24951,g24957,g24958,g24972,g24973,g24974,
    g24975,g24988,g24989,g25002,g25003,g25018,g25019,g25020,g25021,g25038,g25048,g25049,
    g25062,g25172,g25186,I24363,I24364,I24365,g25199,g25200,I24383,I24384,I24385,g25215,
    g25216,g25233,I24414,I24415,I24416,g25236,g25237,g25255,I24438,I24439,I24440,g25258,
    g25268,I24461,I24462,I24463,g25271,g25275,g25293,g25300,g25309,g25334,g25337,g25341,
    g25349,g25381,g25382,g25385,g25389,g25396,g25400,g25425,g25426,g25429,g25432,g25435,
    g25439,g25467,g25470,g25473,g25476,g25492,g25495,g25498,g25514,g25527,g25531,g25532,
    g25537,g25779,g25888,g25895,g25953,g25974,g25984,g25985,g25995,g25996,g26025,g26052,
    g26053,g26208,g26235,I25219,I25220,I25221,g26248,g26255,I25242,I25243,I25244,g26269,
    g26352,g26382,g26666,g26685,g26714,g26745,g26752,g26782,I25845,I25846,I25847,g27141,
    I25907,I25908,I25909,g27223,g27273,g27282,g27295,g27306,g27317,I26049,I26050,I26051,
    g27365,g27377,I26070,I26071,I26072,g27380,I26093,I26094,I26095,g27401,g27463,g27468,
    g27550,g27577,g27582,g27586,g27587,g27593,g27613,g27654,g27670,g27679,g27687,g27693,
    g27705,g27738,I26366,I26367,I26368,g27767,g27775,g27796,I26393,I26394,I26395,g27824,
    g27833,g27854,I26417,I26418,I26419,g27876,g27882,g27903,I26438,I26439,I26440,g27925,
    g27931,g27933,I26459,I26460,I26461,g27955,g28109,g28131,g28167,g28174,g28203,g28206,
    g28207,g28259,g28270,g28271,g28287,g28288,g28298,g28336,g28349,g28363,g28376,g28381,
    g28391,g28395,g28406,g28410,g28421,g28448,g28500,g28504,g28512,g28516,g28522,g28736,
    g28755,g28758,g28765,g28780,g28783,g28786,g28793,g28796,g28820,g28823,g28824,g28827,
    g28830,g28837,g28840,g28843,g28853,g28856,g28857,g28860,g28861,g28864,g28867,g28870,
    g28871,g28874,g28877,g28885,g28888,g28892,g28895,g28896,g28899,g28900,g28903,g28906,
    g28907,g28910,g28911,g28914,g28920,g28923,g28927,g28930,g28931,g28934,g28935,g28938,
    g28942,g28945,g28946,g28949,g28950,g28955,g28958,g28962,g28965,g28966,g28969,g28973,
    g28976,g28977,g28980,g28987,g28990,g28994,g28997,g29001,g29004,g29015,g29018,g29025,
    g29028,g29046,g29049,g29057,g29060,g29082,g29085,g29094,g29097,g29118,g29121,g29131,
    g29134,g29154,g29157,g29186,g29335,g29355,g29540,g29556,g29657,g29660,g29672,g29676,
    g29679,g29694,g29702,g29719,g29722,g29737,g29778,g30573,g30580,g31003,g31009,g31262,
    g31509,I29253,I29254,I29255,g31669,I29261,I29262,I29263,g31671,I29269,I29270,I29271,
    g31706,I29277,I29278,I29279,g31708,I29284,I29285,I29286,g31709,I29295,I29296,I29297,
    g31747,I29302,I29303,I29304,g31748,I29313,I29314,I29315,g31753,g31950,g31971,g31978,
    g31997,g32057,g32072,g33083,g33299,g33306,g33394,g33669,g33679,g33838,g33925,g33930,
    g33933,g34048,I31972,I31973,I31974,g34051,I31983,I31984,I31985,g34056,g34162,g34174,
    I32185,I32186,I32187,g34220,I32202,I32203,I32204,g34227,I32431,I32432,I32433,g34422,
    I32439,I32440,I32441,g34424,I32516,I32517,I32518,g34469,g34545,g34550,I32756,I32757,
    I32758,g34650,g7139,g7142,g7158,g7175,g7192,g7304,g7352,g7499,g7567,g7601,g7661,g7675,
    g7781,g8086,g8131,g8177,g8182,g8720,g8864,g8906,g8933,g8958,g8984,g9015,g9061,g9100,
    g9586,g9602,g9640,g9649,g9664,g9694,g9700,g9755,g9762,g9835,g10123,g10179,g10205,
    g10266,g10281,g10312,g10318,g10338,g10341,g10421,g10488,g10491,g10510,g10555,g10615,
    g10649,g10666,g10671,g10695,g10699,g10709,g10715,g10760,g10793,g10799,g10801,g10803,
    g10808,g10819,g10821,g10831,g10862,g10884,g10893,g10899,g10918,g10922,g11006,g11012,
    g11039,g11107,g11119,g11148,g11171,g11184,g11185,g11191,g11194,g11201,g11203,g11207,
    g11213,g11216,g11217,g11225,g11231,g11232,g11238,g11248,g11252,g11255,g11261,g11270,
    g11273,g11276,g11280,g11283,g11303,g11306,g11309,g11313,g11345,g11346,g11357,g11360,
    g11363,g11384,g11385,g11414,g11415,g11435,g11448,g11469,g11473,g11483,g11493,g11514,
    g11527,g11537,g11563,g11566,g11571,g11584,g11607,g11610,g11618,g11621,g11626,g11653,
    g11658,g11666,g11669,g11692,g11697,g11715,g11729,g11747,g11755,g11763,g11771,g11773,
    g11780,g11797,g11804,g11834,g11846,g11862,g11869,g11885,g11891,g11907,g11913,g11924,
    g11932,g11935,g11940,g11945,g11950,g11954,g11958,g11972,g11976,g11995,g11999,g12002,
    g12017,g12025,g12026,g12029,g12046,g12050,g12059,g12067,g12081,g12085,g12093,g12101,
    g12113,g12117,g12121,g12123,g12126,g12129,g12137,g12146,g12150,g12154,g12160,g12163,
    g12166,g12170,g12173,g12189,g12193,g12198,g12201,g12204,g12208,g12211,g12223,g12226,
    g12228,g12234,g12235,g12246,g12249,g12252,g12256,g12288,g12296,g12297,g12308,g12311,
    g12314,g12318,g12333,g12346,g12347,g12358,g12361,g12364,g12371,g12374,g12377,g12405,
    g12418,g12419,g12432,g12435,g12437,g12443,g12453,g12466,g12467,g12479,g12483,g12486,
    g12492,g12505,g12515,g12540,g12550,g12553,g12558,g12571,g12581,g12591,g12593,g12601,
    g12604,g12609,g12622,g12632,g12645,g12646,g12651,g12659,g12662,g12667,g12680,g12695,
    g12700,g12708,g12711,g12716,g12729,g12739,g12744,g12752,g12755,g12772,g12780,g12785,
    g12798,g12806,g12821,g12824,g12846,g12847,g12848,g12849,g12850,g12851,g12852,g12853,
    g12854,g12855,g12856,g12858,g12970,g12980,g13004,g13005,g13013,g13021,g13031,g13032,
    g13044,g13056,g13076,g13078,g13094,g13110,g13114,g13125,g13129,g13202,g13325,g13326,
    g13335,g13336,g13341,g13342,g13377,g13378,g13480,g13500,g13501,g13512,g13517,g13518,
    g13539,g13568,g13603,g13622,g13631,g13661,g13670,g13698,g13700,g13730,g13765,g13772,
    g13796,g13799,g13806,g13824,g13831,g13852,g13872,g13883,g13908,g13910,g13913,g13919,
    g13937,g13939,g13944,g13946,g13947,g13954,g13959,g13970,g13971,g13989,g13994,g13996,
    g14000,g14001,g14002,g14003,g14027,g14033,g14036,g14037,g14064,g14090,g14091,g14092,
    g14093,g14094,g14121,g14122,g14124,g14145,g14163,g14164,g14165,g14176,g14178,g14181,
    g14188,g14194,g14211,g14212,g14227,g14228,g14247,g14248,g14253,g14271,g14272,g14278,
    g14291,g14306,g14313,g14320,g14334,g14335,g14337,g14339,g14347,g14360,g14361,g14362,
    g14364,g14365,g14367,g14382,g14391,g14392,g14393,g14394,g14395,g14396,g14397,g14399,
    g14411,g14413,g14414,g14415,g14416,g14417,g14418,g14419,g14420,g14425,g14437,g14444,
    g14445,g14446,g14447,g14448,g14449,g14450,g14490,g14497,g14512,g14513,g14514,g14515,
    g14516,g14522,g14529,g14538,g14539,g14540,g14549,g14556,g14568,g14575,g14602,g14611,
    g14640,g14642,g14678,g14679,g14687,g14707,g14712,g14713,g14726,g14731,g14751,g14752,
    g14754,g14767,g14772,g14792,g14793,g14816,g14821,g14867,g14872,g14911,g14914,g14988,
    g15049,g15050,g15051,g15052,g15053,g15054,g15055,g15056,g15057,g15058,g15059,g15060,
    g15061,g15062,g15063,g15064,g15065,g15066,g15067,g15068,g15069,g15070,g15071,g15072,
    g15073,g15074,g15086,g15087,g15088,g15089,g15090,g15091,g15092,g15093,g15094,g15095,
    g15096,g15097,g15098,g15099,g15100,g15101,g15102,g15106,g15120,g15121,g15122,g15123,
    g15126,g15127,g15128,g15129,g15130,g15131,g15132,g15133,g15134,g15135,g15136,g15137,
    g15138,g15139,g15140,g15141,g15142,g15143,g15144,g15145,g15146,g15147,g15148,g15149,
    g15150,g15151,g15152,g15153,g15154,g15155,g15156,g15157,g15158,g15159,g15160,g15161,
    g15162,g15163,g15164,g15165,g15166,g15167,g15168,g15170,g15372,g15508,g15570,g15578,
    g15585,g15594,g15608,g15628,g15647,g15669,g15718,g15724,g15754,g15825,g15992,g16024,
    g16027,g16044,g16066,g16072,g16090,g16183,g16198,g16201,g16209,g16210,g16215,g16219,
    g16220,g16226,g16227,g16231,g16232,g16237,g16242,g16246,g16268,g16272,g16287,g16288,
    g16292,g16313,g16424,g16476,g16479,g16488,g16581,g16646,g17148,g17174,g17175,g17180,
    g17190,g17194,g17198,g17213,g17239,g17284,g17309,g17393,g17420,g17482,g17515,g17619,
    g17625,g17657,g17663,g17694,g17700,g17727,g17954,g19063,g19070,g19140,g19209,g19268,
    g19338,g19388,g19400,g19401,g19402,g19413,g19422,g19430,g19436,g19444,g19453,g19778,
    g19793,g19853,g19873,g19880,g19887,g19890,g19906,g19907,g19919,g19932,g19935,g19951,
    g19953,g19968,g19981,g19984,g19997,g19999,g20000,g20014,g20027,g20149,g20183,g20234,
    g20390,g20717,g20720,g20841,g20854,g20857,g20982,g20995,g20998,g21062,g21127,g21140,
    g21143,g21193,g21206,g21209,g21250,g21256,g21277,g21284,g21389,g21652,g21655,g21658,
    g22190,g22357,g22399,g22400,g22405,g22448,g22450,g22488,g22491,g22513,g22514,g22517,
    g22521,g22522,g22523,g22524,g22535,g22536,g22537,g22539,g22540,g22545,g22654,g22929,
    g22983,g22993,g23024,g23042,g23051,g23052,g23063,g23079,g23108,g23124,g23135,g23204,
    g23208,g23560,g23586,g23602,g23626,g23642,g23662,g23678,g23686,g23695,g23711,g23729,
    g23763,g23835,g23871,g23883,g23918,g23955,g23956,g24018,g24145,g24148,g24383,g24391,
    g24439,g24453,g24494,g24497,g24508,g24514,g24575,g24619,g24631,g24701,g24720,g24751,
    g24766,g24779,g24875,g24953,g24959,g24976,g24990,g25004,g25005,g25022,g25141,g25144,
    g25160,g25175,g25189,g25203,g25247,g25317,g25321,g25407,g25446,g25447,g25501,g25504,
    g25521,g25540,g25769,g25770,g25776,g25777,g25778,g25784,g25785,g25800,g25851,g25887,
    g25932,g25944,g25947,g25948,g25950,g25952,g25954,g25956,g25958,g26098,g26162,g26183,
    g26209,g26212,g26247,g26256,g26267,g26268,g26296,g26297,g26298,g26309,g26314,g26330,
    g26338,g26346,g26515,g26545,g26546,g26573,g26574,g26598,g26603,g26609,g26625,g26628,
    g26645,g26649,g26667,g26686,g26715,g26865,g26872,g26873,g26976,g26993,g27007,g27010,
    g27012,g27027,g27046,g27059,g27063,g27093,g27102,g27337,g27338,g27343,g27344,g27345,
    g27352,g27353,g27354,g27355,g27356,g27364,g27366,g27367,g27368,g27379,g27381,g27382,
    g27400,g27479,g27499,g27511,g27516,g27528,g27629,g27647,g27652,g27659,g27703,g27704,
    g27717,g27720,g27721,g27722,g27731,g27732,g27733,g27734,g27735,g27766,g27768,g27769,
    g27770,g27771,g27772,g27823,g27825,g27826,g27827,g27828,g27829,g27875,g27877,g27878,
    g27879,g27924,g27926,g27927,g27954,g27960,g27966,g27969,g27973,g27982,g28031,g28106,
    g28149,g28340,g28353,g28414,g28425,g28444,g28452,g28457,g28462,g28468,g28469,g28470,
    g28475,g28476,g28480,g28481,g28482,g28483,g28491,g28492,g28493,g28496,g28498,g28509,
    g28510,g28514,g28515,g28519,g28520,g28521,g28529,g28540,g28552,g28568,g28584,g28803,
    g28953,g28981,g28986,g29005,g29006,g29007,g29012,g29032,g29033,g29034,g29035,g29040,
    g29069,g29070,g29071,g29072,g29077,g29104,g29106,g29107,g29108,g29109,g29141,g29142,
    g29144,g29145,g29146,g29164,g29165,g29167,g29173,g29174,g29175,g29179,g29180,g29181,
    g29183,g29184,g29187,g29189,g29191,g29193,g29198,g29200,g29359,g29361,g29370,g29497,
    g29503,g29675,g29705,g29873,g29886,g29889,g29898,g29900,g29903,g29908,g29910,g29915,
    g29916,g29933,g30106,g30117,g30119,g30123,g30129,g30130,g30132,g30134,g30136,g30143,
    g30144,g30146,g30147,g30148,g30150,g30156,g30157,g30159,g30160,g30162,g30169,g30170,
    g30171,g30183,g30240,g30249,g30252,g30260,g30262,g30265,g30271,g30273,g30276,g30280,
    g30282,g30285,g30288,g30290,g30294,g30601,g30613,g30922,g30929,g30934,g31008,g31068,
    g31116,g31117,g31119,g31121,g31126,g31127,g31133,g31134,g31233,g31294,g31318,g31372,
    g31373,g31469,g31476,g31482,g31483,g31491,g31498,g31506,g31507,g31515,g31935,g31942,
    g31965,g31970,g32017,g32212,g32296,g32424,g32455,g32520,g32585,g32650,g32715,g32780,
    g32845,g32910,g33075,g33084,g33085,g33088,g33089,g33090,g33092,g33093,g33094,g33095,
    g33096,g33097,g33098,g33100,g33103,g33107,g33108,g33109,g33112,g33117,g33125,g33128,
    g33129,g33130,g33131,g33132,g33133,g33134,g33135,g33137,g33138,g33139,g33140,g33141,
    g33143,g33144,g33145,g33146,g33147,g33148,g33160,g33161,g33162,g33163,g33174,g33175,
    g33419,g33427,g33432,g33437,g33438,g33439,g33447,g33448,g33449,g33823,g33851,g34067,
    g34354,g34359,g34496,g34703,g34737,g34912;
  dff DFF_1(CK,RST,g72,g24166);
  dff DFF_2(CK,RST,g73,g24167);
  dff DFF_3(CK,RST,g84,g24168);
  dff DFF_4(CK,RST,g90,g24169);
  dff DFF_5(CK,RST,g91,g24170);
  dff DFF_6(CK,RST,g92,g24171);
  dff DFF_7(CK,RST,g99,g24172);
  dff DFF_8(CK,RST,g100,g24173);
  dff DFF_9(CK,RST,g110,g34848);
  dff DFF_10(CK,RST,g112,g34879);
  dff DFF_11(CK,RST,g113,g24174);
  dff DFF_12(CK,RST,g114,g24175);
  dff DFF_13(CK,RST,g115,g24176);
  dff DFF_14(CK,RST,g116,g24177);
  dff DFF_15(CK,RST,g120,g24178);
  dff DFF_16(CK,RST,g124,g24179);
  dff DFF_17(CK,RST,g125,g24180);
  dff DFF_18(CK,RST,g126,g24181);
  dff DFF_19(CK,RST,g127,g24182);
  dff DFF_20(CK,RST,g134,g24183);
  dff DFF_21(CK,RST,g135,g24184);
  dff DFF_22(CK,RST,g44,g24185);
  dff DFF_23(CK,RST,g45,g34990);
  dff DFF_24(CK,RST,g46,g34991);
  dff DFF_25(CK,RST,g47,g34992);
  dff DFF_26(CK,RST,g48,g34993);
  dff DFF_27(CK,RST,g49,g34994);
  dff DFF_28(CK,RST,g50,g34995);
  dff DFF_29(CK,RST,g51,g34996);
  dff DFF_30(CK,RST,g52,g34997);
  dff DFF_31(CK,RST,g53,g24161);
  dff DFF_32(CK,RST,g54,g24162);
  dff DFF_33(CK,RST,g55,g35002);
  dff DFF_34(CK,RST,g56,g24163);
  dff DFF_35(CK,RST,g57,g24164);
  dff DFF_36(CK,RST,g58,g30328);
  dff DFF_37(CK,RST,g63,g34847);
  dff DFF_38(CK,RST,g71,g34786);
  dff DFF_39(CK,RST,g85,g34717);
  dff DFF_40(CK,RST,g93,g34878);
  dff DFF_41(CK,RST,g101,g34787);
  dff DFF_42(CK,RST,g111,g34718);
  dff DFF_43(CK,RST,g43,g34789);
  dff DFF_44(CK,RST,g64,g24165);
  dff DFF_45(CK,RST,g65,g34785);
  dff DFF_46(CK,RST,g70,g18093);
  dff DFF_47(CK,RST,g4507,g30458);
  dff DFF_48(CK,RST,g4459,g34253);
  dff DFF_49(CK,RST,g4369,g26970);
  dff DFF_50(CK,RST,g4473,g34256);
  dff DFF_51(CK,RST,g4462,g34254);
  dff DFF_52(CK,RST,g4581,g26969);
  dff DFF_53(CK,RST,g4467,g34255);
  dff DFF_54(CK,RST,g4474,g10384);
  dff DFF_55(CK,RST,g4477,g26960);
  dff DFF_56(CK,RST,g4480,g31896);
  dff DFF_57(CK,RST,g4495,g33036);
  dff DFF_58(CK,RST,g4498,g33037);
  dff DFF_59(CK,RST,g4501,g33038);
  dff DFF_60(CK,RST,g4504,g33039);
  dff DFF_61(CK,RST,g4512,g33040);
  dff DFF_62(CK,RST,g4521,g26971);
  dff DFF_63(CK,RST,g4527,g28082);
  dff DFF_64(CK,RST,g4515,g26964);
  dff DFF_65(CK,RST,g4519,g33616);
  dff DFF_66(CK,RST,g4520,g6972);
  dff DFF_67(CK,RST,g4483,g4520);
  dff DFF_68(CK,RST,g4486,g26961);
  dff DFF_69(CK,RST,g4489,g26962);
  dff DFF_70(CK,RST,g4492,g26963);
  dff DFF_71(CK,RST,g4537,g34024);
  dff DFF_72(CK,RST,g4423,g4537);
  dff DFF_73(CK,RST,g4540,g31897);
  dff DFF_74(CK,RST,g4543,g33042);
  dff DFF_75(CK,RST,g4567,g33043);
  dff DFF_76(CK,RST,g4546,g33045);
  dff DFF_77(CK,RST,g4549,g33041);
  dff DFF_78(CK,RST,g4552,g33044);
  dff DFF_79(CK,RST,g4570,g33617);
  dff DFF_80(CK,RST,g4571,g6974);
  dff DFF_81(CK,RST,g4555,g4571);
  dff DFF_82(CK,RST,g4558,g26966);
  dff DFF_83(CK,RST,g4561,g26968);
  dff DFF_84(CK,RST,g4564,g26967);
  dff DFF_85(CK,RST,g4534,g34023);
  dff DFF_86(CK,RST,g4420,g26965);
  dff DFF_87(CK,RST,g4438,g26953);
  dff DFF_88(CK,RST,g4449,g26955);
  dff DFF_89(CK,RST,g4443,g4449);
  dff DFF_90(CK,RST,g4446,g26954);
  dff DFF_91(CK,RST,g4452,g4446);
  dff DFF_92(CK,RST,g4434,g26956);
  dff DFF_93(CK,RST,g4430,g26957);
  dff DFF_94(CK,RST,g4427,g26952);
  dff DFF_95(CK,RST,g4375,g26951);
  dff DFF_96(CK,RST,g4414,g26946);
  dff DFF_97(CK,RST,g4411,g4414);
  dff DFF_98(CK,RST,g4408,g26945);
  dff DFF_99(CK,RST,g4405,g4408);
  dff DFF_100(CK,RST,g4401,g26948);
  dff DFF_101(CK,RST,g4388,g26949);
  dff DFF_102(CK,RST,g4382,g26947);
  dff DFF_103(CK,RST,g4417,g31895);
  dff DFF_104(CK,RST,g4392,g26950);
  dff DFF_105(CK,RST,g4456,g25692);
  dff DFF_106(CK,RST,g4455,g26959);
  dff DFF_107(CK,RST,g1,g26958);
  dff DFF_108(CK,RST,g4304,g24281);
  dff DFF_109(CK,RST,g4308,g4304);
  dff DFF_110(CK,RST,g2932,g24282);
  dff DFF_111(CK,RST,g4639,g34025);
  dff DFF_112(CK,RST,g4621,g34460);
  dff DFF_113(CK,RST,g4628,g34457);
  dff DFF_114(CK,RST,g4633,g34458);
  dff DFF_115(CK,RST,g4643,g34259);
  dff DFF_116(CK,RST,g4340,g34459);
  dff DFF_117(CK,RST,g4349,g34257);
  dff DFF_118(CK,RST,g4358,g34258);
  dff DFF_119(CK,RST,g66,g24334);
  dff DFF_120(CK,RST,g4531,g24335);
  dff DFF_121(CK,RST,g4311,g34449);
  dff DFF_122(CK,RST,g4322,g34450);
  dff DFF_123(CK,RST,g4332,g34455);
  dff DFF_124(CK,RST,g4584,g34451);
  dff DFF_125(CK,RST,g4593,g34452);
  dff DFF_126(CK,RST,g4601,g34453);
  dff DFF_127(CK,RST,g4608,g34454);
  dff DFF_128(CK,RST,g4616,g34456);
  dff DFF_129(CK,RST,g4366,g26944);
  dff DFF_130(CK,RST,g4372,g34882);
  dff DFF_131(CK,RST,g4836,g34265);
  dff DFF_132(CK,RST,g4864,g34034);
  dff DFF_133(CK,RST,g4871,g34035);
  dff DFF_134(CK,RST,g4878,g34036);
  dff DFF_135(CK,RST,g4843,g34466);
  dff DFF_136(CK,RST,g4849,g34465);
  dff DFF_137(CK,RST,g4854,g34467);
  dff DFF_138(CK,RST,g4859,g34468);
  dff DFF_139(CK,RST,g4917,g34638);
  dff DFF_140(CK,RST,g4922,g34639);
  dff DFF_141(CK,RST,g4907,g34640);
  dff DFF_142(CK,RST,g4912,g34641);
  dff DFF_143(CK,RST,g4927,g34642);
  dff DFF_144(CK,RST,g4931,g21904);
  dff DFF_145(CK,RST,g4932,g21905);
  dff DFF_146(CK,RST,g4572,g29279);
  dff DFF_147(CK,RST,g4578,g29278);
  dff DFF_148(CK,RST,g4999,g25694);
  dff DFF_149(CK,RST,g5002,g4999);
  dff DFF_150(CK,RST,g5005,g5002);
  dff DFF_151(CK,RST,g5008,g5005);
  dff DFF_152(CK,RST,g4983,g34041);
  dff DFF_153(CK,RST,g4991,g34038);
  dff DFF_154(CK,RST,g4966,g34039);
  dff DFF_155(CK,RST,g4975,g34037);
  dff DFF_156(CK,RST,g4899,g34040);
  dff DFF_157(CK,RST,g4894,g28087);
  dff DFF_158(CK,RST,g4888,g34266);
  dff DFF_159(CK,RST,g4939,g28088);
  dff DFF_160(CK,RST,g4933,g34267);
  dff DFF_161(CK,RST,g4950,g28089);
  dff DFF_162(CK,RST,g4944,g34268);
  dff DFF_163(CK,RST,g4961,g28090);
  dff DFF_164(CK,RST,g4955,g34269);
  dff DFF_165(CK,RST,g4646,g34260);
  dff DFF_166(CK,RST,g4674,g34026);
  dff DFF_167(CK,RST,g4681,g34027);
  dff DFF_168(CK,RST,g4688,g34028);
  dff DFF_169(CK,RST,g4653,g34462);
  dff DFF_170(CK,RST,g4659,g34461);
  dff DFF_171(CK,RST,g4664,g34463);
  dff DFF_172(CK,RST,g4669,g34464);
  dff DFF_173(CK,RST,g4727,g34633);
  dff DFF_174(CK,RST,g4732,g34634);
  dff DFF_175(CK,RST,g4717,g34635);
  dff DFF_176(CK,RST,g4722,g34636);
  dff DFF_177(CK,RST,g4737,g34637);
  dff DFF_178(CK,RST,g4741,g21902);
  dff DFF_179(CK,RST,g4742,g21903);
  dff DFF_180(CK,RST,g59,g29277);
  dff DFF_181(CK,RST,g4575,g29276);
  dff DFF_182(CK,RST,g4809,g25693);
  dff DFF_183(CK,RST,g4812,g4809);
  dff DFF_184(CK,RST,g4815,g4812);
  dff DFF_185(CK,RST,g4818,g4815);
  dff DFF_186(CK,RST,g4793,g34033);
  dff DFF_187(CK,RST,g4801,g34030);
  dff DFF_188(CK,RST,g4776,g34031);
  dff DFF_189(CK,RST,g4785,g34029);
  dff DFF_190(CK,RST,g4709,g34032);
  dff DFF_191(CK,RST,g4704,g28083);
  dff DFF_192(CK,RST,g4698,g34261);
  dff DFF_193(CK,RST,g4749,g28084);
  dff DFF_194(CK,RST,g4743,g34262);
  dff DFF_195(CK,RST,g4760,g28085);
  dff DFF_196(CK,RST,g4754,g34263);
  dff DFF_197(CK,RST,g4771,g28086);
  dff DFF_198(CK,RST,g4765,g34264);
  dff DFF_199(CK,RST,g5313,g24336);
  dff DFF_200(CK,RST,g5290,g5313);
  dff DFF_201(CK,RST,g5320,g5290);
  dff DFF_202(CK,RST,g5276,g5320);
  dff DFF_203(CK,RST,g5283,g5276);
  dff DFF_204(CK,RST,g5308,g5283);
  dff DFF_205(CK,RST,g5327,g5308);
  dff DFF_206(CK,RST,g5331,g5327);
  dff DFF_207(CK,RST,g5335,g5331);
  dff DFF_208(CK,RST,g5339,g5335);
  dff DFF_209(CK,RST,g5343,g24337);
  dff DFF_210(CK,RST,g5348,g24338);
  dff DFF_211(CK,RST,g5352,g24339);
  dff DFF_212(CK,RST,g5357,g33618);
  dff DFF_213(CK,RST,g5297,g33619);
  dff DFF_214(CK,RST,g5101,g25700);
  dff DFF_215(CK,RST,g5109,g5101);
  dff DFF_216(CK,RST,g5062,g25702);
  dff DFF_217(CK,RST,g5105,g25701);
  dff DFF_218(CK,RST,g5112,g5105);
  dff DFF_219(CK,RST,g5022,g25703);
  dff DFF_220(CK,RST,g5016,g31898);
  dff DFF_221(CK,RST,g5029,g31902);
  dff DFF_222(CK,RST,g5033,g31904);
  dff DFF_223(CK,RST,g5037,g31899);
  dff DFF_224(CK,RST,g5041,g31900);
  dff DFF_225(CK,RST,g5046,g31901);
  dff DFF_226(CK,RST,g5052,g31903);
  dff DFF_227(CK,RST,g5057,g33046);
  dff DFF_228(CK,RST,g5069,g28092);
  dff DFF_229(CK,RST,g5073,g28091);
  dff DFF_230(CK,RST,g5077,g25704);
  dff DFF_231(CK,RST,g5080,g25695);
  dff DFF_232(CK,RST,g5084,g25696);
  dff DFF_233(CK,RST,g5092,g25697);
  dff DFF_234(CK,RST,g5097,g25698);
  dff DFF_235(CK,RST,g86,g25699);
  dff DFF_236(CK,RST,g5164,g30459);
  dff DFF_237(CK,RST,g5170,g33047);
  dff DFF_238(CK,RST,g5176,g33048);
  dff DFF_239(CK,RST,g5180,g33049);
  dff DFF_240(CK,RST,g5188,g33050);
  dff DFF_241(CK,RST,g5196,g30460);
  dff DFF_242(CK,RST,g5224,g30464);
  dff DFF_243(CK,RST,g5240,g30468);
  dff DFF_244(CK,RST,g5256,g30472);
  dff DFF_245(CK,RST,g5204,g30476);
  dff DFF_246(CK,RST,g5200,g30461);
  dff DFF_247(CK,RST,g5228,g30465);
  dff DFF_248(CK,RST,g5244,g30469);
  dff DFF_249(CK,RST,g5260,g30473);
  dff DFF_250(CK,RST,g5212,g30477);
  dff DFF_251(CK,RST,g5208,g30462);
  dff DFF_252(CK,RST,g5232,g30466);
  dff DFF_253(CK,RST,g5248,g30470);
  dff DFF_254(CK,RST,g5264,g30474);
  dff DFF_255(CK,RST,g5220,g30478);
  dff DFF_256(CK,RST,g5216,g30463);
  dff DFF_257(CK,RST,g5236,g30467);
  dff DFF_258(CK,RST,g5252,g30471);
  dff DFF_259(CK,RST,g5268,g30475);
  dff DFF_260(CK,RST,g5272,g30479);
  dff DFF_261(CK,RST,g128,g28093);
  dff DFF_262(CK,RST,g5156,g29285);
  dff DFF_263(CK,RST,g5120,g25708);
  dff DFF_264(CK,RST,g5115,g29280);
  dff DFF_265(CK,RST,g5124,g29281);
  dff DFF_266(CK,RST,g5128,g25705);
  dff DFF_267(CK,RST,g5134,g29282);
  dff DFF_268(CK,RST,g5138,g29283);
  dff DFF_269(CK,RST,g5142,g29284);
  dff DFF_270(CK,RST,g5148,g25706);
  dff DFF_271(CK,RST,g5152,g25707);
  dff DFF_272(CK,RST,g5160,g34643);
  dff DFF_273(CK,RST,g5659,g24340);
  dff DFF_274(CK,RST,g5637,g5659);
  dff DFF_275(CK,RST,g5666,g5637);
  dff DFF_276(CK,RST,g5623,g5666);
  dff DFF_277(CK,RST,g5630,g5623);
  dff DFF_278(CK,RST,g5654,g5630);
  dff DFF_279(CK,RST,g5673,g5654);
  dff DFF_280(CK,RST,g5677,g5673);
  dff DFF_281(CK,RST,g5681,g5677);
  dff DFF_282(CK,RST,g5685,g5681);
  dff DFF_283(CK,RST,g5689,g24341);
  dff DFF_284(CK,RST,g5694,g24342);
  dff DFF_285(CK,RST,g5698,g24343);
  dff DFF_286(CK,RST,g5703,g33620);
  dff DFF_287(CK,RST,g5644,g33621);
  dff DFF_288(CK,RST,g5448,g25714);
  dff DFF_289(CK,RST,g5456,g5448);
  dff DFF_290(CK,RST,g5406,g25716);
  dff DFF_291(CK,RST,g5452,g25715);
  dff DFF_292(CK,RST,g5459,g5452);
  dff DFF_293(CK,RST,g5366,g25717);
  dff DFF_294(CK,RST,g5360,g31905);
  dff DFF_295(CK,RST,g5373,g31909);
  dff DFF_296(CK,RST,g5377,g31911);
  dff DFF_297(CK,RST,g5381,g31906);
  dff DFF_298(CK,RST,g5385,g31907);
  dff DFF_299(CK,RST,g5390,g31908);
  dff DFF_300(CK,RST,g5396,g31910);
  dff DFF_301(CK,RST,g5401,g33051);
  dff DFF_302(CK,RST,g5413,g28095);
  dff DFF_303(CK,RST,g5417,g28094);
  dff DFF_304(CK,RST,g5421,g25718);
  dff DFF_305(CK,RST,g5424,g25709);
  dff DFF_306(CK,RST,g5428,g25710);
  dff DFF_307(CK,RST,g5436,g25711);
  dff DFF_308(CK,RST,g5441,g25712);
  dff DFF_309(CK,RST,g5445,g25713);
  dff DFF_310(CK,RST,g5511,g30480);
  dff DFF_311(CK,RST,g5517,g33052);
  dff DFF_312(CK,RST,g5523,g33053);
  dff DFF_313(CK,RST,g5527,g33054);
  dff DFF_314(CK,RST,g5535,g33055);
  dff DFF_315(CK,RST,g5543,g30481);
  dff DFF_316(CK,RST,g5571,g30485);
  dff DFF_317(CK,RST,g5587,g30489);
  dff DFF_318(CK,RST,g5603,g30493);
  dff DFF_319(CK,RST,g5551,g30497);
  dff DFF_320(CK,RST,g5547,g30482);
  dff DFF_321(CK,RST,g5575,g30486);
  dff DFF_322(CK,RST,g5591,g30490);
  dff DFF_323(CK,RST,g5607,g30494);
  dff DFF_324(CK,RST,g5559,g30498);
  dff DFF_325(CK,RST,g5555,g30483);
  dff DFF_326(CK,RST,g5579,g30487);
  dff DFF_327(CK,RST,g5595,g30491);
  dff DFF_328(CK,RST,g5611,g30495);
  dff DFF_329(CK,RST,g5567,g30499);
  dff DFF_330(CK,RST,g5563,g30484);
  dff DFF_331(CK,RST,g5583,g30488);
  dff DFF_332(CK,RST,g5599,g30492);
  dff DFF_333(CK,RST,g5615,g30496);
  dff DFF_334(CK,RST,g5619,g30500);
  dff DFF_335(CK,RST,g4821,g28096);
  dff DFF_336(CK,RST,g5503,g29291);
  dff DFF_337(CK,RST,g5467,g25722);
  dff DFF_338(CK,RST,g5462,g29286);
  dff DFF_339(CK,RST,g5471,g29287);
  dff DFF_340(CK,RST,g5475,g25719);
  dff DFF_341(CK,RST,g5481,g29288);
  dff DFF_342(CK,RST,g5485,g29289);
  dff DFF_343(CK,RST,g5489,g29290);
  dff DFF_344(CK,RST,g5495,g25720);
  dff DFF_345(CK,RST,g5499,g25721);
  dff DFF_346(CK,RST,g5507,g34644);
  dff DFF_347(CK,RST,g6005,g24344);
  dff DFF_348(CK,RST,g5983,g6005);
  dff DFF_349(CK,RST,g6012,g5983);
  dff DFF_350(CK,RST,g5969,g6012);
  dff DFF_351(CK,RST,g5976,g5969);
  dff DFF_352(CK,RST,g6000,g5976);
  dff DFF_353(CK,RST,g6019,g6000);
  dff DFF_354(CK,RST,g6023,g6019);
  dff DFF_355(CK,RST,g6027,g6023);
  dff DFF_356(CK,RST,g6031,g6027);
  dff DFF_357(CK,RST,g6035,g24345);
  dff DFF_358(CK,RST,g6040,g24346);
  dff DFF_359(CK,RST,g6044,g24347);
  dff DFF_360(CK,RST,g6049,g33622);
  dff DFF_361(CK,RST,g5990,g33623);
  dff DFF_362(CK,RST,g5794,g25728);
  dff DFF_363(CK,RST,g5802,g5794);
  dff DFF_364(CK,RST,g5752,g25730);
  dff DFF_365(CK,RST,g5798,g25729);
  dff DFF_366(CK,RST,g5805,g5798);
  dff DFF_367(CK,RST,g5712,g25731);
  dff DFF_368(CK,RST,g5706,g31912);
  dff DFF_369(CK,RST,g5719,g31916);
  dff DFF_370(CK,RST,g5723,g31918);
  dff DFF_371(CK,RST,g5727,g31913);
  dff DFF_372(CK,RST,g5731,g31914);
  dff DFF_373(CK,RST,g5736,g31915);
  dff DFF_374(CK,RST,g5742,g31917);
  dff DFF_375(CK,RST,g5747,g33056);
  dff DFF_376(CK,RST,g5759,g28098);
  dff DFF_377(CK,RST,g5763,g28097);
  dff DFF_378(CK,RST,g5767,g25732);
  dff DFF_379(CK,RST,g5770,g25723);
  dff DFF_380(CK,RST,g5774,g25724);
  dff DFF_381(CK,RST,g5782,g25725);
  dff DFF_382(CK,RST,g5787,g25726);
  dff DFF_383(CK,RST,g5791,g25727);
  dff DFF_384(CK,RST,g5857,g30501);
  dff DFF_385(CK,RST,g5863,g33057);
  dff DFF_386(CK,RST,g5869,g33058);
  dff DFF_387(CK,RST,g5873,g33059);
  dff DFF_388(CK,RST,g5881,g33060);
  dff DFF_389(CK,RST,g5889,g30502);
  dff DFF_390(CK,RST,g5917,g30506);
  dff DFF_391(CK,RST,g5933,g30510);
  dff DFF_392(CK,RST,g5949,g30514);
  dff DFF_393(CK,RST,g5897,g30518);
  dff DFF_394(CK,RST,g5893,g30503);
  dff DFF_395(CK,RST,g5921,g30507);
  dff DFF_396(CK,RST,g5937,g30511);
  dff DFF_397(CK,RST,g5953,g30515);
  dff DFF_398(CK,RST,g5905,g30519);
  dff DFF_399(CK,RST,g5901,g30504);
  dff DFF_400(CK,RST,g5925,g30508);
  dff DFF_401(CK,RST,g5941,g30512);
  dff DFF_402(CK,RST,g5957,g30516);
  dff DFF_403(CK,RST,g5913,g30520);
  dff DFF_404(CK,RST,g5909,g30505);
  dff DFF_405(CK,RST,g5929,g30509);
  dff DFF_406(CK,RST,g5945,g30513);
  dff DFF_407(CK,RST,g5961,g30517);
  dff DFF_408(CK,RST,g5965,g30521);
  dff DFF_409(CK,RST,g4831,g28099);
  dff DFF_410(CK,RST,g5849,g29297);
  dff DFF_411(CK,RST,g5813,g25736);
  dff DFF_412(CK,RST,g5808,g29292);
  dff DFF_413(CK,RST,g5817,g29293);
  dff DFF_414(CK,RST,g5821,g25733);
  dff DFF_415(CK,RST,g5827,g29294);
  dff DFF_416(CK,RST,g5831,g29295);
  dff DFF_417(CK,RST,g5835,g29296);
  dff DFF_418(CK,RST,g5841,g25734);
  dff DFF_419(CK,RST,g5845,g25735);
  dff DFF_420(CK,RST,g5853,g34645);
  dff DFF_421(CK,RST,g6351,g24348);
  dff DFF_422(CK,RST,g6329,g6351);
  dff DFF_423(CK,RST,g6358,g6329);
  dff DFF_424(CK,RST,g6315,g6358);
  dff DFF_425(CK,RST,g6322,g6315);
  dff DFF_426(CK,RST,g6346,g6322);
  dff DFF_427(CK,RST,g6365,g6346);
  dff DFF_428(CK,RST,g6369,g6365);
  dff DFF_429(CK,RST,g6373,g6369);
  dff DFF_430(CK,RST,g6377,g6373);
  dff DFF_431(CK,RST,g6381,g24349);
  dff DFF_432(CK,RST,g6386,g24350);
  dff DFF_433(CK,RST,g6390,g24351);
  dff DFF_434(CK,RST,g6395,g33624);
  dff DFF_435(CK,RST,g6336,g33625);
  dff DFF_436(CK,RST,g6140,g25742);
  dff DFF_437(CK,RST,g6148,g6140);
  dff DFF_438(CK,RST,g6098,g25744);
  dff DFF_439(CK,RST,g6144,g25743);
  dff DFF_440(CK,RST,g6151,g6144);
  dff DFF_441(CK,RST,g6058,g25745);
  dff DFF_442(CK,RST,g6052,g31919);
  dff DFF_443(CK,RST,g6065,g31923);
  dff DFF_444(CK,RST,g6069,g31925);
  dff DFF_445(CK,RST,g6073,g31920);
  dff DFF_446(CK,RST,g6077,g31921);
  dff DFF_447(CK,RST,g6082,g31922);
  dff DFF_448(CK,RST,g6088,g31924);
  dff DFF_449(CK,RST,g6093,g33061);
  dff DFF_450(CK,RST,g6105,g28101);
  dff DFF_451(CK,RST,g6109,g28100);
  dff DFF_452(CK,RST,g6113,g25746);
  dff DFF_453(CK,RST,g6116,g25737);
  dff DFF_454(CK,RST,g6120,g25738);
  dff DFF_455(CK,RST,g6128,g25739);
  dff DFF_456(CK,RST,g6133,g25740);
  dff DFF_457(CK,RST,g6137,g25741);
  dff DFF_458(CK,RST,g6203,g30522);
  dff DFF_459(CK,RST,g6209,g33062);
  dff DFF_460(CK,RST,g6215,g33063);
  dff DFF_461(CK,RST,g6219,g33064);
  dff DFF_462(CK,RST,g6227,g33065);
  dff DFF_463(CK,RST,g6235,g30523);
  dff DFF_464(CK,RST,g6263,g30527);
  dff DFF_465(CK,RST,g6279,g30531);
  dff DFF_466(CK,RST,g6295,g30535);
  dff DFF_467(CK,RST,g6243,g30539);
  dff DFF_468(CK,RST,g6239,g30524);
  dff DFF_469(CK,RST,g6267,g30528);
  dff DFF_470(CK,RST,g6283,g30532);
  dff DFF_471(CK,RST,g6299,g30536);
  dff DFF_472(CK,RST,g6251,g30540);
  dff DFF_473(CK,RST,g6247,g30525);
  dff DFF_474(CK,RST,g6271,g30529);
  dff DFF_475(CK,RST,g6287,g30533);
  dff DFF_476(CK,RST,g6303,g30537);
  dff DFF_477(CK,RST,g6259,g30541);
  dff DFF_478(CK,RST,g6255,g30526);
  dff DFF_479(CK,RST,g6275,g30530);
  dff DFF_480(CK,RST,g6291,g30534);
  dff DFF_481(CK,RST,g6307,g30538);
  dff DFF_482(CK,RST,g6311,g30542);
  dff DFF_483(CK,RST,g4826,g28102);
  dff DFF_484(CK,RST,g6195,g29303);
  dff DFF_485(CK,RST,g6159,g25750);
  dff DFF_486(CK,RST,g6154,g29298);
  dff DFF_487(CK,RST,g6163,g29299);
  dff DFF_488(CK,RST,g6167,g25747);
  dff DFF_489(CK,RST,g6173,g29300);
  dff DFF_490(CK,RST,g6177,g29301);
  dff DFF_491(CK,RST,g6181,g29302);
  dff DFF_492(CK,RST,g6187,g25748);
  dff DFF_493(CK,RST,g6191,g25749);
  dff DFF_494(CK,RST,g6199,g34646);
  dff DFF_495(CK,RST,g6697,g24352);
  dff DFF_496(CK,RST,g6675,g6697);
  dff DFF_497(CK,RST,g6704,g6675);
  dff DFF_498(CK,RST,g6661,g6704);
  dff DFF_499(CK,RST,g6668,g6661);
  dff DFF_500(CK,RST,g6692,g6668);
  dff DFF_501(CK,RST,g6711,g6692);
  dff DFF_502(CK,RST,g6715,g6711);
  dff DFF_503(CK,RST,g6719,g6715);
  dff DFF_504(CK,RST,g6723,g6719);
  dff DFF_505(CK,RST,g6727,g24353);
  dff DFF_506(CK,RST,g6732,g24354);
  dff DFF_507(CK,RST,g6736,g24355);
  dff DFF_508(CK,RST,g6741,g33626);
  dff DFF_509(CK,RST,g6682,g33627);
  dff DFF_510(CK,RST,g6486,g25756);
  dff DFF_511(CK,RST,g6494,g6486);
  dff DFF_512(CK,RST,g6444,g25758);
  dff DFF_513(CK,RST,g6490,g25757);
  dff DFF_514(CK,RST,g6497,g6490);
  dff DFF_515(CK,RST,g6404,g25759);
  dff DFF_516(CK,RST,g6398,g31926);
  dff DFF_517(CK,RST,g6411,g31930);
  dff DFF_518(CK,RST,g6415,g31932);
  dff DFF_519(CK,RST,g6419,g31927);
  dff DFF_520(CK,RST,g6423,g31928);
  dff DFF_521(CK,RST,g6428,g31929);
  dff DFF_522(CK,RST,g6434,g31931);
  dff DFF_523(CK,RST,g6439,g33066);
  dff DFF_524(CK,RST,g6451,g28104);
  dff DFF_525(CK,RST,g6455,g28103);
  dff DFF_526(CK,RST,g6459,g25760);
  dff DFF_527(CK,RST,g6462,g25751);
  dff DFF_528(CK,RST,g6466,g25752);
  dff DFF_529(CK,RST,g6474,g25753);
  dff DFF_530(CK,RST,g6479,g25754);
  dff DFF_531(CK,RST,g6483,g25755);
  dff DFF_532(CK,RST,g6549,g30543);
  dff DFF_533(CK,RST,g6555,g33067);
  dff DFF_534(CK,RST,g6561,g33068);
  dff DFF_535(CK,RST,g6565,g33069);
  dff DFF_536(CK,RST,g6573,g33070);
  dff DFF_537(CK,RST,g6581,g30544);
  dff DFF_538(CK,RST,g6609,g30548);
  dff DFF_539(CK,RST,g6625,g30552);
  dff DFF_540(CK,RST,g6641,g30556);
  dff DFF_541(CK,RST,g6589,g30560);
  dff DFF_542(CK,RST,g6585,g30545);
  dff DFF_543(CK,RST,g6613,g30549);
  dff DFF_544(CK,RST,g6629,g30553);
  dff DFF_545(CK,RST,g6645,g30557);
  dff DFF_546(CK,RST,g6597,g30561);
  dff DFF_547(CK,RST,g6593,g30546);
  dff DFF_548(CK,RST,g6617,g30550);
  dff DFF_549(CK,RST,g6633,g30554);
  dff DFF_550(CK,RST,g6649,g30558);
  dff DFF_551(CK,RST,g6605,g30562);
  dff DFF_552(CK,RST,g6601,g30547);
  dff DFF_553(CK,RST,g6621,g30551);
  dff DFF_554(CK,RST,g6637,g30555);
  dff DFF_555(CK,RST,g6653,g30559);
  dff DFF_556(CK,RST,g6657,g30563);
  dff DFF_557(CK,RST,g5011,g28105);
  dff DFF_558(CK,RST,g6541,g29309);
  dff DFF_559(CK,RST,g6505,g25764);
  dff DFF_560(CK,RST,g6500,g29304);
  dff DFF_561(CK,RST,g6509,g29305);
  dff DFF_562(CK,RST,g6513,g25761);
  dff DFF_563(CK,RST,g6519,g29306);
  dff DFF_564(CK,RST,g6523,g29307);
  dff DFF_565(CK,RST,g6527,g29308);
  dff DFF_566(CK,RST,g6533,g25762);
  dff DFF_567(CK,RST,g6537,g25763);
  dff DFF_568(CK,RST,g6545,g34647);
  dff DFF_569(CK,RST,g3303,g24267);
  dff DFF_570(CK,RST,g3281,g3303);
  dff DFF_571(CK,RST,g3310,g3281);
  dff DFF_572(CK,RST,g3267,g3310);
  dff DFF_573(CK,RST,g3274,g3267);
  dff DFF_574(CK,RST,g3298,g3274);
  dff DFF_575(CK,RST,g3317,g3298);
  dff DFF_576(CK,RST,g3321,g3317);
  dff DFF_577(CK,RST,g3325,g3321);
  dff DFF_578(CK,RST,g3329,g3325);
  dff DFF_579(CK,RST,g3338,g24268);
  dff DFF_580(CK,RST,g3343,g24269);
  dff DFF_581(CK,RST,g3347,g24270);
  dff DFF_582(CK,RST,g3352,g33609);
  dff DFF_583(CK,RST,g3288,g33610);
  dff DFF_584(CK,RST,g3092,g25648);
  dff DFF_585(CK,RST,g3100,g3092);
  dff DFF_586(CK,RST,g3050,g25650);
  dff DFF_587(CK,RST,g3096,g25649);
  dff DFF_588(CK,RST,g3103,g3096);
  dff DFF_589(CK,RST,g3010,g25651);
  dff DFF_590(CK,RST,g3004,g31873);
  dff DFF_591(CK,RST,g3017,g31877);
  dff DFF_592(CK,RST,g3021,g31879);
  dff DFF_593(CK,RST,g3025,g31874);
  dff DFF_594(CK,RST,g3029,g31875);
  dff DFF_595(CK,RST,g3034,g31876);
  dff DFF_596(CK,RST,g3040,g31878);
  dff DFF_597(CK,RST,g3045,g33020);
  dff DFF_598(CK,RST,g3057,g28062);
  dff DFF_599(CK,RST,g3061,g28061);
  dff DFF_600(CK,RST,g3065,g25652);
  dff DFF_601(CK,RST,g3068,g25643);
  dff DFF_602(CK,RST,g3072,g25644);
  dff DFF_603(CK,RST,g3080,g25645);
  dff DFF_604(CK,RST,g3085,g25646);
  dff DFF_605(CK,RST,g3089,g25647);
  dff DFF_606(CK,RST,g3155,g30393);
  dff DFF_607(CK,RST,g3161,g33021);
  dff DFF_608(CK,RST,g3167,g33022);
  dff DFF_609(CK,RST,g3171,g33023);
  dff DFF_610(CK,RST,g3179,g33024);
  dff DFF_611(CK,RST,g3187,g30394);
  dff DFF_612(CK,RST,g3215,g30398);
  dff DFF_613(CK,RST,g3231,g30402);
  dff DFF_614(CK,RST,g3247,g30406);
  dff DFF_615(CK,RST,g3195,g30410);
  dff DFF_616(CK,RST,g3191,g30395);
  dff DFF_617(CK,RST,g3219,g30399);
  dff DFF_618(CK,RST,g3235,g30403);
  dff DFF_619(CK,RST,g3251,g30407);
  dff DFF_620(CK,RST,g3203,g30411);
  dff DFF_621(CK,RST,g3199,g30396);
  dff DFF_622(CK,RST,g3223,g30400);
  dff DFF_623(CK,RST,g3239,g30404);
  dff DFF_624(CK,RST,g3255,g30408);
  dff DFF_625(CK,RST,g3211,g30412);
  dff DFF_626(CK,RST,g3207,g30397);
  dff DFF_627(CK,RST,g3227,g30401);
  dff DFF_628(CK,RST,g3243,g30405);
  dff DFF_629(CK,RST,g3259,g30409);
  dff DFF_630(CK,RST,g3263,g30413);
  dff DFF_631(CK,RST,g3333,g28063);
  dff DFF_632(CK,RST,g3147,g29262);
  dff DFF_633(CK,RST,g3111,g25656);
  dff DFF_634(CK,RST,g3106,g29257);
  dff DFF_635(CK,RST,g3115,g29258);
  dff DFF_636(CK,RST,g3119,g25653);
  dff DFF_637(CK,RST,g3125,g29259);
  dff DFF_638(CK,RST,g3129,g29260);
  dff DFF_639(CK,RST,g3133,g29261);
  dff DFF_640(CK,RST,g3139,g25654);
  dff DFF_641(CK,RST,g3143,g25655);
  dff DFF_642(CK,RST,g3151,g34625);
  dff DFF_643(CK,RST,g3654,g24271);
  dff DFF_644(CK,RST,g3632,g3654);
  dff DFF_645(CK,RST,g3661,g3632);
  dff DFF_646(CK,RST,g3618,g3661);
  dff DFF_647(CK,RST,g3625,g3618);
  dff DFF_648(CK,RST,g3649,g3625);
  dff DFF_649(CK,RST,g3668,g3649);
  dff DFF_650(CK,RST,g3672,g3668);
  dff DFF_651(CK,RST,g3676,g3672);
  dff DFF_652(CK,RST,g3680,g3676);
  dff DFF_653(CK,RST,g3689,g24272);
  dff DFF_654(CK,RST,g3694,g24273);
  dff DFF_655(CK,RST,g3698,g24274);
  dff DFF_656(CK,RST,g3703,g33611);
  dff DFF_657(CK,RST,g3639,g33612);
  dff DFF_658(CK,RST,g3443,g25662);
  dff DFF_659(CK,RST,g3451,g3443);
  dff DFF_660(CK,RST,g3401,g25664);
  dff DFF_661(CK,RST,g3447,g25663);
  dff DFF_662(CK,RST,g3454,g3447);
  dff DFF_663(CK,RST,g3361,g25665);
  dff DFF_664(CK,RST,g3355,g31880);
  dff DFF_665(CK,RST,g3368,g31884);
  dff DFF_666(CK,RST,g3372,g31886);
  dff DFF_667(CK,RST,g3376,g31881);
  dff DFF_668(CK,RST,g3380,g31882);
  dff DFF_669(CK,RST,g3385,g31883);
  dff DFF_670(CK,RST,g3391,g31885);
  dff DFF_671(CK,RST,g3396,g33025);
  dff DFF_672(CK,RST,g3408,g28065);
  dff DFF_673(CK,RST,g3412,g28064);
  dff DFF_674(CK,RST,g3416,g25666);
  dff DFF_675(CK,RST,g3419,g25657);
  dff DFF_676(CK,RST,g3423,g25658);
  dff DFF_677(CK,RST,g3431,g25659);
  dff DFF_678(CK,RST,g3436,g25660);
  dff DFF_679(CK,RST,g3440,g25661);
  dff DFF_680(CK,RST,g3506,g30414);
  dff DFF_681(CK,RST,g3512,g33026);
  dff DFF_682(CK,RST,g3518,g33027);
  dff DFF_683(CK,RST,g3522,g33028);
  dff DFF_684(CK,RST,g3530,g33029);
  dff DFF_685(CK,RST,g3538,g30415);
  dff DFF_686(CK,RST,g3566,g30419);
  dff DFF_687(CK,RST,g3582,g30423);
  dff DFF_688(CK,RST,g3598,g30427);
  dff DFF_689(CK,RST,g3546,g30431);
  dff DFF_690(CK,RST,g3542,g30416);
  dff DFF_691(CK,RST,g3570,g30420);
  dff DFF_692(CK,RST,g3586,g30424);
  dff DFF_693(CK,RST,g3602,g30428);
  dff DFF_694(CK,RST,g3554,g30432);
  dff DFF_695(CK,RST,g3550,g30417);
  dff DFF_696(CK,RST,g3574,g30421);
  dff DFF_697(CK,RST,g3590,g30425);
  dff DFF_698(CK,RST,g3606,g30429);
  dff DFF_699(CK,RST,g3562,g30433);
  dff DFF_700(CK,RST,g3558,g30418);
  dff DFF_701(CK,RST,g3578,g30422);
  dff DFF_702(CK,RST,g3594,g30426);
  dff DFF_703(CK,RST,g3610,g30430);
  dff DFF_704(CK,RST,g3614,g30434);
  dff DFF_705(CK,RST,g3684,g28066);
  dff DFF_706(CK,RST,g3498,g29268);
  dff DFF_707(CK,RST,g3462,g25670);
  dff DFF_708(CK,RST,g3457,g29263);
  dff DFF_709(CK,RST,g3466,g29264);
  dff DFF_710(CK,RST,g3470,g25667);
  dff DFF_711(CK,RST,g3476,g29265);
  dff DFF_712(CK,RST,g3480,g29266);
  dff DFF_713(CK,RST,g3484,g29267);
  dff DFF_714(CK,RST,g3490,g25668);
  dff DFF_715(CK,RST,g3494,g25669);
  dff DFF_716(CK,RST,g3502,g34626);
  dff DFF_717(CK,RST,g4005,g24275);
  dff DFF_718(CK,RST,g3983,g4005);
  dff DFF_719(CK,RST,g4012,g3983);
  dff DFF_720(CK,RST,g3969,g4012);
  dff DFF_721(CK,RST,g3976,g3969);
  dff DFF_722(CK,RST,g4000,g3976);
  dff DFF_723(CK,RST,g4019,g4000);
  dff DFF_724(CK,RST,g4023,g4019);
  dff DFF_725(CK,RST,g4027,g4023);
  dff DFF_726(CK,RST,g4031,g4027);
  dff DFF_727(CK,RST,g4040,g24276);
  dff DFF_728(CK,RST,g4045,g24277);
  dff DFF_729(CK,RST,g4049,g24278);
  dff DFF_730(CK,RST,g4054,g33613);
  dff DFF_731(CK,RST,g3990,g33614);
  dff DFF_732(CK,RST,g3794,g25676);
  dff DFF_733(CK,RST,g3802,g3794);
  dff DFF_734(CK,RST,g3752,g25678);
  dff DFF_735(CK,RST,g3798,g25677);
  dff DFF_736(CK,RST,g3805,g3798);
  dff DFF_737(CK,RST,g3712,g25679);
  dff DFF_738(CK,RST,g3706,g31887);
  dff DFF_739(CK,RST,g3719,g31891);
  dff DFF_740(CK,RST,g3723,g31893);
  dff DFF_741(CK,RST,g3727,g31888);
  dff DFF_742(CK,RST,g3731,g31889);
  dff DFF_743(CK,RST,g3736,g31890);
  dff DFF_744(CK,RST,g3742,g31892);
  dff DFF_745(CK,RST,g3747,g33030);
  dff DFF_746(CK,RST,g3759,g28068);
  dff DFF_747(CK,RST,g3763,g28067);
  dff DFF_748(CK,RST,g3767,g25680);
  dff DFF_749(CK,RST,g3770,g25671);
  dff DFF_750(CK,RST,g3774,g25672);
  dff DFF_751(CK,RST,g3782,g25673);
  dff DFF_752(CK,RST,g3787,g25674);
  dff DFF_753(CK,RST,g3791,g25675);
  dff DFF_754(CK,RST,g3857,g30435);
  dff DFF_755(CK,RST,g3863,g33031);
  dff DFF_756(CK,RST,g3869,g33032);
  dff DFF_757(CK,RST,g3873,g33033);
  dff DFF_758(CK,RST,g3881,g33034);
  dff DFF_759(CK,RST,g3889,g30436);
  dff DFF_760(CK,RST,g3917,g30440);
  dff DFF_761(CK,RST,g3933,g30444);
  dff DFF_762(CK,RST,g3949,g30448);
  dff DFF_763(CK,RST,g3897,g30452);
  dff DFF_764(CK,RST,g3893,g30437);
  dff DFF_765(CK,RST,g3921,g30441);
  dff DFF_766(CK,RST,g3937,g30445);
  dff DFF_767(CK,RST,g3953,g30449);
  dff DFF_768(CK,RST,g3905,g30453);
  dff DFF_769(CK,RST,g3901,g30438);
  dff DFF_770(CK,RST,g3925,g30442);
  dff DFF_771(CK,RST,g3941,g30446);
  dff DFF_772(CK,RST,g3957,g30450);
  dff DFF_773(CK,RST,g3913,g30454);
  dff DFF_774(CK,RST,g3909,g30439);
  dff DFF_775(CK,RST,g3929,g30443);
  dff DFF_776(CK,RST,g3945,g30447);
  dff DFF_777(CK,RST,g3961,g30451);
  dff DFF_778(CK,RST,g3965,g30455);
  dff DFF_779(CK,RST,g4035,g28069);
  dff DFF_780(CK,RST,g3849,g29274);
  dff DFF_781(CK,RST,g3813,g25684);
  dff DFF_782(CK,RST,g3808,g29269);
  dff DFF_783(CK,RST,g3817,g29270);
  dff DFF_784(CK,RST,g3821,g25681);
  dff DFF_785(CK,RST,g3827,g29271);
  dff DFF_786(CK,RST,g3831,g29272);
  dff DFF_787(CK,RST,g3835,g29273);
  dff DFF_788(CK,RST,g3841,g25682);
  dff DFF_789(CK,RST,g3845,g25683);
  dff DFF_790(CK,RST,g3853,g34627);
  dff DFF_791(CK,RST,g4165,g28079);
  dff DFF_792(CK,RST,g4169,g28080);
  dff DFF_793(CK,RST,g4125,g28081);
  dff DFF_794(CK,RST,g4072,g25691);
  dff DFF_795(CK,RST,g4064,g25685);
  dff DFF_796(CK,RST,g4057,g25686);
  dff DFF_797(CK,RST,g4141,g25687);
  dff DFF_798(CK,RST,g4082,g26938);
  dff DFF_799(CK,RST,g4076,g28070);
  dff DFF_800(CK,RST,g4087,g29275);
  dff DFF_801(CK,RST,g4093,g30456);
  dff DFF_802(CK,RST,g4098,g31894);
  dff DFF_803(CK,RST,g4108,g33035);
  dff DFF_804(CK,RST,g4104,g33615);
  dff DFF_805(CK,RST,g4145,g26939);
  dff DFF_806(CK,RST,g4112,g28071);
  dff DFF_807(CK,RST,g4116,g28072);
  dff DFF_808(CK,RST,g4119,g28073);
  dff DFF_809(CK,RST,g4122,g28074);
  dff DFF_810(CK,RST,g4153,g30457);
  dff DFF_811(CK,RST,g4164,g26940);
  dff DFF_812(CK,RST,g4129,g28075);
  dff DFF_813(CK,RST,g4132,g28076);
  dff DFF_814(CK,RST,g4135,g28077);
  dff DFF_815(CK,RST,g4138,g28078);
  dff DFF_816(CK,RST,g4172,g34733);
  dff DFF_817(CK,RST,g4176,g34734);
  dff DFF_818(CK,RST,g4146,g34628);
  dff DFF_819(CK,RST,g4157,g34629);
  dff DFF_820(CK,RST,g4258,g21893);
  dff DFF_821(CK,RST,g4264,g21894);
  dff DFF_822(CK,RST,g4269,g21895);
  dff DFF_823(CK,RST,g4273,g24280);
  dff DFF_824(CK,RST,g4239,g21892);
  dff DFF_825(CK,RST,g4294,g21900);
  dff DFF_826(CK,RST,g4297,g4294);
  dff DFF_827(CK,RST,g4300,g34735);
  dff DFF_828(CK,RST,g4253,g34630);
  dff DFF_829(CK,RST,g4249,g34631);
  dff DFF_830(CK,RST,g4245,g34632);
  dff DFF_831(CK,RST,g4277,g21896);
  dff DFF_832(CK,RST,g4281,g4277);
  dff DFF_833(CK,RST,g4284,g21897);
  dff DFF_834(CK,RST,g4287,g21898);
  dff DFF_835(CK,RST,g4291,g4287);
  dff DFF_836(CK,RST,g2946,g21899);
  dff DFF_837(CK,RST,g4191,g21901);
  dff DFF_838(CK,RST,g4188,g4191);
  dff DFF_839(CK,RST,g4194,g4188);
  dff DFF_840(CK,RST,g4197,g4194);
  dff DFF_841(CK,RST,g4200,g4197);
  dff DFF_842(CK,RST,g4204,g4200);
  dff DFF_843(CK,RST,g4207,g4204);
  dff DFF_844(CK,RST,g4210,g4207);
  dff DFF_845(CK,RST,g4180,g4210);
  dff DFF_846(CK,RST,g4185,g21891);
  dff DFF_847(CK,RST,g4213,g4185);
  dff DFF_848(CK,RST,g4216,g4213);
  dff DFF_849(CK,RST,g4219,g4216);
  dff DFF_850(CK,RST,g4222,g4219);
  dff DFF_851(CK,RST,g4226,g4222);
  dff DFF_852(CK,RST,g4229,g4226);
  dff DFF_853(CK,RST,g4232,g4229);
  dff DFF_854(CK,RST,g4235,g4232);
  dff DFF_855(CK,RST,g4242,g24279);
  dff DFF_856(CK,RST,g305,g26880);
  dff DFF_857(CK,RST,g311,g26881);
  dff DFF_858(CK,RST,g336,g26886);
  dff DFF_859(CK,RST,g324,g26887);
  dff DFF_860(CK,RST,g316,g26883);
  dff DFF_861(CK,RST,g319,g26882);
  dff DFF_862(CK,RST,g329,g26885);
  dff DFF_863(CK,RST,g333,g26884);
  dff DFF_864(CK,RST,g344,g26890);
  dff DFF_865(CK,RST,g347,g344);
  dff DFF_866(CK,RST,g351,g26891);
  dff DFF_867(CK,RST,g355,g26892);
  dff DFF_868(CK,RST,g74,g26893);
  dff DFF_869(CK,RST,g106,g26889);
  dff DFF_870(CK,RST,g341,g26888);
  dff DFF_871(CK,RST,g637,g24212);
  dff DFF_872(CK,RST,g640,g637);
  dff DFF_873(CK,RST,g559,g640);
  dff DFF_874(CK,RST,g562,g25613);
  dff DFF_875(CK,RST,g568,g26895);
  dff DFF_876(CK,RST,g572,g28045);
  dff DFF_877(CK,RST,g586,g29224);
  dff DFF_878(CK,RST,g577,g30334);
  dff DFF_879(CK,RST,g582,g31866);
  dff DFF_880(CK,RST,g590,g32978);
  dff DFF_881(CK,RST,g595,g33538);
  dff DFF_882(CK,RST,g599,g33964);
  dff DFF_883(CK,RST,g604,g34251);
  dff DFF_884(CK,RST,g608,g34438);
  dff DFF_885(CK,RST,g613,g34599);
  dff DFF_886(CK,RST,g617,g34724);
  dff DFF_887(CK,RST,g622,g34790);
  dff DFF_888(CK,RST,g626,g34849);
  dff DFF_889(CK,RST,g632,g34880);
  dff DFF_890(CK,RST,g859,g26900);
  dff DFF_891(CK,RST,g869,g859);
  dff DFF_892(CK,RST,g875,g869);
  dff DFF_893(CK,RST,g878,g875);
  dff DFF_894(CK,RST,g881,g878);
  dff DFF_895(CK,RST,g884,g881);
  dff DFF_896(CK,RST,g887,g884);
  dff DFF_897(CK,RST,g872,g887);
  dff DFF_898(CK,RST,g225,g26901);
  dff DFF_899(CK,RST,g255,g26902);
  dff DFF_900(CK,RST,g232,g26903);
  dff DFF_901(CK,RST,g262,g26904);
  dff DFF_902(CK,RST,g239,g26905);
  dff DFF_903(CK,RST,g269,g26906);
  dff DFF_904(CK,RST,g246,g26907);
  dff DFF_905(CK,RST,g446,g26908);
  dff DFF_906(CK,RST,g890,g34440);
  dff DFF_907(CK,RST,g862,g26909);
  dff DFF_908(CK,RST,g896,g26910);
  dff DFF_909(CK,RST,g901,g25620);
  dff DFF_910(CK,RST,g391,g26911);
  dff DFF_911(CK,RST,g365,g25595);
  dff DFF_912(CK,RST,g358,g365);
  dff DFF_913(CK,RST,g370,g25597);
  dff DFF_914(CK,RST,g376,g25596);
  dff DFF_915(CK,RST,g385,g25598);
  dff DFF_916(CK,RST,g203,g25599);
  dff DFF_917(CK,RST,g854,g32980);
  dff DFF_918(CK,RST,g847,g24216);
  dff DFF_919(CK,RST,g703,g24214);
  dff DFF_920(CK,RST,g837,g24215);
  dff DFF_921(CK,RST,g843,g25619);
  dff DFF_922(CK,RST,g812,g26898);
  dff DFF_923(CK,RST,g817,g25617);
  dff DFF_924(CK,RST,g832,g25618);
  dff DFF_925(CK,RST,g822,g26899);
  dff DFF_926(CK,RST,g827,g28055);
  dff DFF_927(CK,RST,g723,g29229);
  dff DFF_928(CK,RST,g645,g28046);
  dff DFF_929(CK,RST,g681,g28047);
  dff DFF_930(CK,RST,g699,g28053);
  dff DFF_931(CK,RST,g650,g28049);
  dff DFF_932(CK,RST,g655,g28050);
  dff DFF_933(CK,RST,g718,g28051);
  dff DFF_934(CK,RST,g661,g28052);
  dff DFF_935(CK,RST,g728,g28054);
  dff DFF_936(CK,RST,g79,g26896);
  dff DFF_937(CK,RST,g691,g28048);
  dff DFF_938(CK,RST,g686,g25614);
  dff DFF_939(CK,RST,g667,g25615);
  dff DFF_940(CK,RST,g671,g29225);
  dff DFF_941(CK,RST,g676,g29226);
  dff DFF_942(CK,RST,g714,g29227);
  dff DFF_943(CK,RST,g499,g25609);
  dff DFF_944(CK,RST,g504,g25610);
  dff DFF_945(CK,RST,g513,g25611);
  dff DFF_946(CK,RST,g518,g25612);
  dff DFF_947(CK,RST,g528,g26894);
  dff DFF_948(CK,RST,g482,g28044);
  dff DFF_949(CK,RST,g490,g29223);
  dff DFF_950(CK,RST,g417,g24209);
  dff DFF_951(CK,RST,g411,g29222);
  dff DFF_952(CK,RST,g424,g24202);
  dff DFF_953(CK,RST,g475,g24208);
  dff DFF_954(CK,RST,g441,g24207);
  dff DFF_955(CK,RST,g437,g24206);
  dff DFF_956(CK,RST,g433,g24205);
  dff DFF_957(CK,RST,g429,g24204);
  dff DFF_958(CK,RST,g401,g24203);
  dff DFF_959(CK,RST,g392,g24200);
  dff DFF_960(CK,RST,g405,g24201);
  dff DFF_961(CK,RST,g182,g25602);
  dff DFF_962(CK,RST,g174,g25601);
  dff DFF_963(CK,RST,g168,g25600);
  dff DFF_964(CK,RST,g460,g25605);
  dff DFF_965(CK,RST,g452,g25604);
  dff DFF_966(CK,RST,g457,g25603);
  dff DFF_967(CK,RST,g471,g25608);
  dff DFF_968(CK,RST,g464,g25607);
  dff DFF_969(CK,RST,g468,g25606);
  dff DFF_970(CK,RST,g479,g24210);
  dff DFF_971(CK,RST,g102,g33962);
  dff DFF_972(CK,RST,g496,g33963);
  dff DFF_973(CK,RST,g732,g25616);
  dff DFF_974(CK,RST,g753,g26897);
  dff DFF_975(CK,RST,g799,g24213);
  dff DFF_976(CK,RST,g802,g799);
  dff DFF_977(CK,RST,g736,g802);
  dff DFF_978(CK,RST,g739,g29228);
  dff DFF_979(CK,RST,g744,g30335);
  dff DFF_980(CK,RST,g749,g31867);
  dff DFF_981(CK,RST,g758,g32979);
  dff DFF_982(CK,RST,g763,g33539);
  dff DFF_983(CK,RST,g767,g33965);
  dff DFF_984(CK,RST,g772,g34252);
  dff DFF_985(CK,RST,g776,g34439);
  dff DFF_986(CK,RST,g781,g34600);
  dff DFF_987(CK,RST,g785,g34725);
  dff DFF_988(CK,RST,g790,g34791);
  dff DFF_989(CK,RST,g794,g34850);
  dff DFF_990(CK,RST,g807,g34881);
  dff DFF_991(CK,RST,g554,g34911);
  dff DFF_992(CK,RST,g538,g34719);
  dff DFF_993(CK,RST,g546,g34722);
  dff DFF_994(CK,RST,g542,g24211);
  dff DFF_995(CK,RST,g534,g34723);
  dff DFF_996(CK,RST,g550,g34720);
  dff DFF_997(CK,RST,g136,g34598);
  dff DFF_998(CK,RST,g199,g34721);
  dff DFF_999(CK,RST,g278,g25594);
  dff DFF_1000(CK,RST,g283,g28043);
  dff DFF_1001(CK,RST,g287,g31865);
  dff DFF_1002(CK,RST,g291,g32977);
  dff DFF_1003(CK,RST,g294,g33535);
  dff DFF_1004(CK,RST,g298,g33961);
  dff DFF_1005(CK,RST,g142,g34250);
  dff DFF_1006(CK,RST,g146,g30333);
  dff DFF_1007(CK,RST,g164,g31864);
  dff DFF_1008(CK,RST,g150,g32976);
  dff DFF_1009(CK,RST,g153,g33534);
  dff DFF_1010(CK,RST,g157,g33960);
  dff DFF_1011(CK,RST,g160,g34249);
  dff DFF_1012(CK,RST,g301,g33536);
  dff DFF_1013(CK,RST,g222,g33537);
  dff DFF_1014(CK,RST,g194,g25592);
  dff DFF_1015(CK,RST,g191,g194);
  dff DFF_1016(CK,RST,g209,g25593);
  dff DFF_1017(CK,RST,g215,g25591);
  dff DFF_1018(CK,RST,g218,g215);
  dff DFF_1019(CK,RST,g1249,g24247);
  dff DFF_1020(CK,RST,g1266,g25630);
  dff DFF_1021(CK,RST,g1280,g26919);
  dff DFF_1022(CK,RST,g1252,g28058);
  dff DFF_1023(CK,RST,g1256,g29235);
  dff DFF_1024(CK,RST,g1259,g30342);
  dff DFF_1025(CK,RST,g1263,g31870);
  dff DFF_1026(CK,RST,g1270,g32984);
  dff DFF_1027(CK,RST,g1274,g33542);
  dff DFF_1028(CK,RST,g1277,g32985);
  dff DFF_1029(CK,RST,g1418,g24254);
  dff DFF_1030(CK,RST,g1422,g1418);
  dff DFF_1031(CK,RST,g1426,g1422);
  dff DFF_1032(CK,RST,g1430,g1426);
  dff DFF_1033(CK,RST,g1548,g24260);
  dff DFF_1034(CK,RST,g1564,g24262);
  dff DFF_1035(CK,RST,g1559,g25638);
  dff DFF_1036(CK,RST,g1554,g25637);
  dff DFF_1037(CK,RST,g1570,g24258);
  dff DFF_1038(CK,RST,g1585,g1570);
  dff DFF_1039(CK,RST,g1589,g24261);
  dff DFF_1040(CK,RST,g1576,g24255);
  dff DFF_1041(CK,RST,g1579,g1576);
  dff DFF_1042(CK,RST,g1339,g24259);
  dff DFF_1043(CK,RST,g1500,g24256);
  dff DFF_1044(CK,RST,g1582,g1500);
  dff DFF_1045(CK,RST,g1333,g1582);
  dff DFF_1046(CK,RST,g1399,g24257);
  dff DFF_1047(CK,RST,g1459,g1399);
  dff DFF_1048(CK,RST,g1322,g1459);
  dff DFF_1049(CK,RST,g1514,g30344);
  dff DFF_1050(CK,RST,g1526,g30345);
  dff DFF_1051(CK,RST,g1521,g24252);
  dff DFF_1052(CK,RST,g1306,g25636);
  dff DFF_1053(CK,RST,g1532,g24253);
  dff DFF_1054(CK,RST,g1536,g26925);
  dff DFF_1055(CK,RST,g1542,g30346);
  dff DFF_1056(CK,RST,g1413,g30347);
  dff DFF_1057(CK,RST,g1395,g25634);
  dff DFF_1058(CK,RST,g1404,g26921);
  dff DFF_1059(CK,RST,g1319,g24248);
  dff DFF_1060(CK,RST,g1312,g25631);
  dff DFF_1061(CK,RST,g1351,g25632);
  dff DFF_1062(CK,RST,g1345,g28059);
  dff DFF_1063(CK,RST,g1361,g30343);
  dff DFF_1064(CK,RST,g1367,g31871);
  dff DFF_1065(CK,RST,g1373,g32986);
  dff DFF_1066(CK,RST,g1379,g33543);
  dff DFF_1067(CK,RST,g1384,g25633);
  dff DFF_1068(CK,RST,g1389,g26920);
  dff DFF_1069(CK,RST,g1489,g24249);
  dff DFF_1070(CK,RST,g1495,g24250);
  dff DFF_1071(CK,RST,g1442,g24251);
  dff DFF_1072(CK,RST,g1437,g29236);
  dff DFF_1073(CK,RST,g1478,g26924);
  dff DFF_1074(CK,RST,g1454,g29239);
  dff DFF_1075(CK,RST,g1448,g26922);
  dff DFF_1076(CK,RST,g1467,g29237);
  dff DFF_1077(CK,RST,g1472,g26923);
  dff DFF_1078(CK,RST,g1484,g29238);
  dff DFF_1079(CK,RST,g1300,g25635);
  dff DFF_1080(CK,RST,g1291,g34602);
  dff DFF_1081(CK,RST,g1296,g34729);
  dff DFF_1082(CK,RST,g1283,g34730);
  dff DFF_1083(CK,RST,g1287,g34731);
  dff DFF_1084(CK,RST,g1311,g21724);
  dff DFF_1085(CK,RST,g929,g21725);
  dff DFF_1086(CK,RST,g904,g24231);
  dff DFF_1087(CK,RST,g921,g25621);
  dff DFF_1088(CK,RST,g936,g26912);
  dff DFF_1089(CK,RST,g907,g28056);
  dff DFF_1090(CK,RST,g911,g29230);
  dff DFF_1091(CK,RST,g914,g30336);
  dff DFF_1092(CK,RST,g918,g31868);
  dff DFF_1093(CK,RST,g925,g32981);
  dff DFF_1094(CK,RST,g930,g33540);
  dff DFF_1095(CK,RST,g933,g32982);
  dff DFF_1096(CK,RST,g1075,g24238);
  dff DFF_1097(CK,RST,g1079,g1075);
  dff DFF_1098(CK,RST,g1083,g1079);
  dff DFF_1099(CK,RST,g1087,g1083);
  dff DFF_1100(CK,RST,g1205,g24244);
  dff DFF_1101(CK,RST,g1221,g24246);
  dff DFF_1102(CK,RST,g1216,g25629);
  dff DFF_1103(CK,RST,g1211,g25628);
  dff DFF_1104(CK,RST,g1227,g24242);
  dff DFF_1105(CK,RST,g1242,g1227);
  dff DFF_1106(CK,RST,g1246,g24245);
  dff DFF_1107(CK,RST,g1233,g24239);
  dff DFF_1108(CK,RST,g1236,g1233);
  dff DFF_1109(CK,RST,g996,g24243);
  dff DFF_1110(CK,RST,g1157,g24240);
  dff DFF_1111(CK,RST,g1239,g1157);
  dff DFF_1112(CK,RST,g990,g1239);
  dff DFF_1113(CK,RST,g1056,g24241);
  dff DFF_1114(CK,RST,g1116,g1056);
  dff DFF_1115(CK,RST,g979,g1116);
  dff DFF_1116(CK,RST,g1171,g30338);
  dff DFF_1117(CK,RST,g1183,g30339);
  dff DFF_1118(CK,RST,g1178,g24236);
  dff DFF_1119(CK,RST,g962,g25627);
  dff DFF_1120(CK,RST,g1189,g24237);
  dff DFF_1121(CK,RST,g1193,g26918);
  dff DFF_1122(CK,RST,g1199,g30340);
  dff DFF_1123(CK,RST,g1070,g30341);
  dff DFF_1124(CK,RST,g1052,g25625);
  dff DFF_1125(CK,RST,g1061,g26914);
  dff DFF_1126(CK,RST,g976,g24232);
  dff DFF_1127(CK,RST,g969,g25622);
  dff DFF_1128(CK,RST,g1008,g25623);
  dff DFF_1129(CK,RST,g1002,g28057);
  dff DFF_1130(CK,RST,g1018,g30337);
  dff DFF_1131(CK,RST,g1024,g31869);
  dff DFF_1132(CK,RST,g1030,g32983);
  dff DFF_1133(CK,RST,g1036,g33541);
  dff DFF_1134(CK,RST,g1041,g25624);
  dff DFF_1135(CK,RST,g1046,g26913);
  dff DFF_1136(CK,RST,g1146,g24233);
  dff DFF_1137(CK,RST,g1152,g24234);
  dff DFF_1138(CK,RST,g1099,g24235);
  dff DFF_1139(CK,RST,g1094,g29231);
  dff DFF_1140(CK,RST,g1135,g26917);
  dff DFF_1141(CK,RST,g1111,g29234);
  dff DFF_1142(CK,RST,g1105,g26915);
  dff DFF_1143(CK,RST,g1124,g29232);
  dff DFF_1144(CK,RST,g1129,g26916);
  dff DFF_1145(CK,RST,g1141,g29233);
  dff DFF_1146(CK,RST,g956,g25626);
  dff DFF_1147(CK,RST,g947,g34601);
  dff DFF_1148(CK,RST,g952,g34726);
  dff DFF_1149(CK,RST,g939,g34727);
  dff DFF_1150(CK,RST,g943,g34728);
  dff DFF_1151(CK,RST,g967,g21722);
  dff DFF_1152(CK,RST,g968,g21723);
  dff DFF_1153(CK,RST,g1592,g33544);
  dff DFF_1154(CK,RST,g1644,g33551);
  dff DFF_1155(CK,RST,g1636,g33545);
  dff DFF_1156(CK,RST,g1668,g33546);
  dff DFF_1157(CK,RST,g1682,g33971);
  dff DFF_1158(CK,RST,g1687,g33547);
  dff DFF_1159(CK,RST,g1604,g33972);
  dff DFF_1160(CK,RST,g1600,g33966);
  dff DFF_1161(CK,RST,g1608,g33967);
  dff DFF_1162(CK,RST,g1620,g33970);
  dff DFF_1163(CK,RST,g1616,g33969);
  dff DFF_1164(CK,RST,g1612,g33968);
  dff DFF_1165(CK,RST,g1632,g30348);
  dff DFF_1166(CK,RST,g1624,g32987);
  dff DFF_1167(CK,RST,g1648,g32988);
  dff DFF_1168(CK,RST,g1664,g32990);
  dff DFF_1169(CK,RST,g1657,g32989);
  dff DFF_1170(CK,RST,g1677,g29240);
  dff DFF_1171(CK,RST,g1691,g29241);
  dff DFF_1172(CK,RST,g1696,g30349);
  dff DFF_1173(CK,RST,g1700,g30350);
  dff DFF_1174(CK,RST,g1706,g33548);
  dff DFF_1175(CK,RST,g1710,g33549);
  dff DFF_1176(CK,RST,g1714,g33550);
  dff DFF_1177(CK,RST,g1720,g30351);
  dff DFF_1178(CK,RST,g1724,g30352);
  dff DFF_1179(CK,RST,g1728,g33552);
  dff DFF_1180(CK,RST,g1779,g33559);
  dff DFF_1181(CK,RST,g1772,g33553);
  dff DFF_1182(CK,RST,g1802,g33554);
  dff DFF_1183(CK,RST,g1816,g33978);
  dff DFF_1184(CK,RST,g1821,g33555);
  dff DFF_1185(CK,RST,g1740,g33979);
  dff DFF_1186(CK,RST,g1736,g33973);
  dff DFF_1187(CK,RST,g1744,g33974);
  dff DFF_1188(CK,RST,g1756,g33977);
  dff DFF_1189(CK,RST,g1752,g33976);
  dff DFF_1190(CK,RST,g1748,g33975);
  dff DFF_1191(CK,RST,g1768,g30353);
  dff DFF_1192(CK,RST,g1760,g32991);
  dff DFF_1193(CK,RST,g1783,g32992);
  dff DFF_1194(CK,RST,g1798,g32994);
  dff DFF_1195(CK,RST,g1792,g32993);
  dff DFF_1196(CK,RST,g1811,g29242);
  dff DFF_1197(CK,RST,g1825,g29243);
  dff DFF_1198(CK,RST,g1830,g30354);
  dff DFF_1199(CK,RST,g1834,g30355);
  dff DFF_1200(CK,RST,g1840,g33556);
  dff DFF_1201(CK,RST,g1844,g33557);
  dff DFF_1202(CK,RST,g1848,g33558);
  dff DFF_1203(CK,RST,g1854,g30356);
  dff DFF_1204(CK,RST,g1858,g30357);
  dff DFF_1205(CK,RST,g1862,g33560);
  dff DFF_1206(CK,RST,g1913,g33567);
  dff DFF_1207(CK,RST,g1906,g33561);
  dff DFF_1208(CK,RST,g1936,g33562);
  dff DFF_1209(CK,RST,g1950,g33985);
  dff DFF_1210(CK,RST,g1955,g33563);
  dff DFF_1211(CK,RST,g1874,g33986);
  dff DFF_1212(CK,RST,g1870,g33980);
  dff DFF_1213(CK,RST,g1878,g33981);
  dff DFF_1214(CK,RST,g1890,g33984);
  dff DFF_1215(CK,RST,g1886,g33983);
  dff DFF_1216(CK,RST,g1882,g33982);
  dff DFF_1217(CK,RST,g1902,g30358);
  dff DFF_1218(CK,RST,g1894,g32995);
  dff DFF_1219(CK,RST,g1917,g32996);
  dff DFF_1220(CK,RST,g1932,g32998);
  dff DFF_1221(CK,RST,g1926,g32997);
  dff DFF_1222(CK,RST,g1945,g29244);
  dff DFF_1223(CK,RST,g1959,g29245);
  dff DFF_1224(CK,RST,g1964,g30359);
  dff DFF_1225(CK,RST,g1968,g30360);
  dff DFF_1226(CK,RST,g1974,g33564);
  dff DFF_1227(CK,RST,g1978,g33565);
  dff DFF_1228(CK,RST,g1982,g33566);
  dff DFF_1229(CK,RST,g1988,g30361);
  dff DFF_1230(CK,RST,g1992,g30362);
  dff DFF_1231(CK,RST,g1996,g33568);
  dff DFF_1232(CK,RST,g2047,g33575);
  dff DFF_1233(CK,RST,g2040,g33569);
  dff DFF_1234(CK,RST,g2070,g33570);
  dff DFF_1235(CK,RST,g2084,g33992);
  dff DFF_1236(CK,RST,g2089,g33571);
  dff DFF_1237(CK,RST,g2008,g33993);
  dff DFF_1238(CK,RST,g2004,g33987);
  dff DFF_1239(CK,RST,g2012,g33988);
  dff DFF_1240(CK,RST,g2024,g33991);
  dff DFF_1241(CK,RST,g2020,g33990);
  dff DFF_1242(CK,RST,g2016,g33989);
  dff DFF_1243(CK,RST,g2036,g30363);
  dff DFF_1244(CK,RST,g2028,g32999);
  dff DFF_1245(CK,RST,g2051,g33000);
  dff DFF_1246(CK,RST,g2066,g33002);
  dff DFF_1247(CK,RST,g2060,g33001);
  dff DFF_1248(CK,RST,g2079,g29246);
  dff DFF_1249(CK,RST,g2093,g29247);
  dff DFF_1250(CK,RST,g2098,g30364);
  dff DFF_1251(CK,RST,g2102,g30365);
  dff DFF_1252(CK,RST,g2108,g33572);
  dff DFF_1253(CK,RST,g2112,g33573);
  dff DFF_1254(CK,RST,g2116,g33574);
  dff DFF_1255(CK,RST,g2122,g30366);
  dff DFF_1256(CK,RST,g2126,g30367);
  dff DFF_1257(CK,RST,g2130,g34603);
  dff DFF_1258(CK,RST,g2138,g34604);
  dff DFF_1259(CK,RST,g2145,g34605);
  dff DFF_1260(CK,RST,g2151,g18421);
  dff DFF_1261(CK,RST,g2152,g18422);
  dff DFF_1262(CK,RST,g2153,g33576);
  dff DFF_1263(CK,RST,g2204,g33583);
  dff DFF_1264(CK,RST,g2197,g33577);
  dff DFF_1265(CK,RST,g2227,g33578);
  dff DFF_1266(CK,RST,g2241,g33999);
  dff DFF_1267(CK,RST,g2246,g33579);
  dff DFF_1268(CK,RST,g2165,g34000);
  dff DFF_1269(CK,RST,g2161,g33994);
  dff DFF_1270(CK,RST,g2169,g33995);
  dff DFF_1271(CK,RST,g2181,g33998);
  dff DFF_1272(CK,RST,g2177,g33997);
  dff DFF_1273(CK,RST,g2173,g33996);
  dff DFF_1274(CK,RST,g2193,g30368);
  dff DFF_1275(CK,RST,g2185,g33003);
  dff DFF_1276(CK,RST,g2208,g33004);
  dff DFF_1277(CK,RST,g2223,g33006);
  dff DFF_1278(CK,RST,g2217,g33005);
  dff DFF_1279(CK,RST,g2236,g29248);
  dff DFF_1280(CK,RST,g2250,g29249);
  dff DFF_1281(CK,RST,g2255,g30369);
  dff DFF_1282(CK,RST,g2259,g30370);
  dff DFF_1283(CK,RST,g2265,g33580);
  dff DFF_1284(CK,RST,g2269,g33581);
  dff DFF_1285(CK,RST,g2273,g33582);
  dff DFF_1286(CK,RST,g2279,g30371);
  dff DFF_1287(CK,RST,g2283,g30372);
  dff DFF_1288(CK,RST,g2287,g33584);
  dff DFF_1289(CK,RST,g2338,g33591);
  dff DFF_1290(CK,RST,g2331,g33585);
  dff DFF_1291(CK,RST,g2361,g33586);
  dff DFF_1292(CK,RST,g2375,g34006);
  dff DFF_1293(CK,RST,g2380,g33587);
  dff DFF_1294(CK,RST,g2299,g34007);
  dff DFF_1295(CK,RST,g2295,g34001);
  dff DFF_1296(CK,RST,g2303,g34002);
  dff DFF_1297(CK,RST,g2315,g34005);
  dff DFF_1298(CK,RST,g2311,g34004);
  dff DFF_1299(CK,RST,g2307,g34003);
  dff DFF_1300(CK,RST,g2327,g30373);
  dff DFF_1301(CK,RST,g2319,g33007);
  dff DFF_1302(CK,RST,g2342,g33008);
  dff DFF_1303(CK,RST,g2357,g33010);
  dff DFF_1304(CK,RST,g2351,g33009);
  dff DFF_1305(CK,RST,g2370,g29250);
  dff DFF_1306(CK,RST,g2384,g29251);
  dff DFF_1307(CK,RST,g2389,g30374);
  dff DFF_1308(CK,RST,g2393,g30375);
  dff DFF_1309(CK,RST,g2399,g33588);
  dff DFF_1310(CK,RST,g2403,g33589);
  dff DFF_1311(CK,RST,g2407,g33590);
  dff DFF_1312(CK,RST,g2413,g30376);
  dff DFF_1313(CK,RST,g2417,g30377);
  dff DFF_1314(CK,RST,g2421,g33592);
  dff DFF_1315(CK,RST,g2472,g33599);
  dff DFF_1316(CK,RST,g2465,g33593);
  dff DFF_1317(CK,RST,g2495,g33594);
  dff DFF_1318(CK,RST,g2509,g34013);
  dff DFF_1319(CK,RST,g2514,g33595);
  dff DFF_1320(CK,RST,g2433,g34014);
  dff DFF_1321(CK,RST,g2429,g34008);
  dff DFF_1322(CK,RST,g2437,g34009);
  dff DFF_1323(CK,RST,g2449,g34012);
  dff DFF_1324(CK,RST,g2445,g34011);
  dff DFF_1325(CK,RST,g2441,g34010);
  dff DFF_1326(CK,RST,g2461,g30378);
  dff DFF_1327(CK,RST,g2453,g33011);
  dff DFF_1328(CK,RST,g2476,g33012);
  dff DFF_1329(CK,RST,g2491,g33014);
  dff DFF_1330(CK,RST,g2485,g33013);
  dff DFF_1331(CK,RST,g2504,g29252);
  dff DFF_1332(CK,RST,g2518,g29253);
  dff DFF_1333(CK,RST,g2523,g30379);
  dff DFF_1334(CK,RST,g2527,g30380);
  dff DFF_1335(CK,RST,g2533,g33596);
  dff DFF_1336(CK,RST,g2537,g33597);
  dff DFF_1337(CK,RST,g2541,g33598);
  dff DFF_1338(CK,RST,g2547,g30381);
  dff DFF_1339(CK,RST,g2551,g30382);
  dff DFF_1340(CK,RST,g2555,g33600);
  dff DFF_1341(CK,RST,g2606,g33607);
  dff DFF_1342(CK,RST,g2599,g33601);
  dff DFF_1343(CK,RST,g2629,g33602);
  dff DFF_1344(CK,RST,g2643,g34020);
  dff DFF_1345(CK,RST,g2648,g33603);
  dff DFF_1346(CK,RST,g2567,g34021);
  dff DFF_1347(CK,RST,g2563,g34015);
  dff DFF_1348(CK,RST,g2571,g34016);
  dff DFF_1349(CK,RST,g2583,g34019);
  dff DFF_1350(CK,RST,g2579,g34018);
  dff DFF_1351(CK,RST,g2575,g34017);
  dff DFF_1352(CK,RST,g2595,g30383);
  dff DFF_1353(CK,RST,g2587,g33015);
  dff DFF_1354(CK,RST,g2610,g33016);
  dff DFF_1355(CK,RST,g2625,g33018);
  dff DFF_1356(CK,RST,g2619,g33017);
  dff DFF_1357(CK,RST,g2638,g29254);
  dff DFF_1358(CK,RST,g2652,g29255);
  dff DFF_1359(CK,RST,g2657,g30384);
  dff DFF_1360(CK,RST,g2661,g30385);
  dff DFF_1361(CK,RST,g2667,g33604);
  dff DFF_1362(CK,RST,g2671,g33605);
  dff DFF_1363(CK,RST,g2675,g33606);
  dff DFF_1364(CK,RST,g2681,g30386);
  dff DFF_1365(CK,RST,g2685,g30387);
  dff DFF_1366(CK,RST,g2689,g34606);
  dff DFF_1367(CK,RST,g2697,g34607);
  dff DFF_1368(CK,RST,g2704,g34608);
  dff DFF_1369(CK,RST,g2710,g18527);
  dff DFF_1370(CK,RST,g2711,g18528);
  dff DFF_1371(CK,RST,g2837,g26935);
  dff DFF_1372(CK,RST,g2841,g26936);
  dff DFF_1373(CK,RST,g2712,g26937);
  dff DFF_1374(CK,RST,g2715,g24263);
  dff DFF_1375(CK,RST,g2719,g25639);
  dff DFF_1376(CK,RST,g2724,g26926);
  dff DFF_1377(CK,RST,g2729,g28060);
  dff DFF_1378(CK,RST,g2735,g29256);
  dff DFF_1379(CK,RST,g2741,g30388);
  dff DFF_1380(CK,RST,g2748,g31872);
  dff DFF_1381(CK,RST,g2756,g33019);
  dff DFF_1382(CK,RST,g2759,g33608);
  dff DFF_1383(CK,RST,g2763,g34022);
  dff DFF_1384(CK,RST,g2767,g26927);
  dff DFF_1385(CK,RST,g2779,g26928);
  dff DFF_1386(CK,RST,g2791,g26929);
  dff DFF_1387(CK,RST,g2795,g26930);
  dff DFF_1388(CK,RST,g2787,g34444);
  dff DFF_1389(CK,RST,g2783,g34442);
  dff DFF_1390(CK,RST,g2775,g34443);
  dff DFF_1391(CK,RST,g2771,g34441);
  dff DFF_1392(CK,RST,g2831,g30391);
  dff DFF_1393(CK,RST,g121,g30389);
  dff DFF_1394(CK,RST,g2799,g26931);
  dff DFF_1395(CK,RST,g2811,g26932);
  dff DFF_1396(CK,RST,g2823,g26933);
  dff DFF_1397(CK,RST,g2827,g26934);
  dff DFF_1398(CK,RST,g2819,g34448);
  dff DFF_1399(CK,RST,g2815,g34446);
  dff DFF_1400(CK,RST,g2807,g34447);
  dff DFF_1401(CK,RST,g2803,g34445);
  dff DFF_1402(CK,RST,g2834,g30392);
  dff DFF_1403(CK,RST,g117,g30390);
  dff DFF_1404(CK,RST,g2999,g34805);
  dff DFF_1405(CK,RST,g2994,g34732);
  dff DFF_1406(CK,RST,g2988,g34624);
  dff DFF_1407(CK,RST,g2868,g34616);
  dff DFF_1408(CK,RST,g2873,g34615);
  dff DFF_1409(CK,RST,g2890,g34799);
  dff DFF_1410(CK,RST,g2844,g34609);
  dff DFF_1411(CK,RST,g2852,g34610);
  dff DFF_1412(CK,RST,g2860,g34611);
  dff DFF_1413(CK,RST,g2894,g34612);
  dff DFF_1414(CK,RST,g37,g34613);
  dff DFF_1415(CK,RST,g94,g34614);
  dff DFF_1416(CK,RST,g2848,g34792);
  dff DFF_1417(CK,RST,g2856,g34793);
  dff DFF_1418(CK,RST,g2864,g34794);
  dff DFF_1419(CK,RST,g2898,g34795);
  dff DFF_1420(CK,RST,g2882,g34796);
  dff DFF_1421(CK,RST,g2878,g34797);
  dff DFF_1422(CK,RST,g2886,g34798);
  dff DFF_1423(CK,RST,g2980,g34800);
  dff DFF_1424(CK,RST,g2984,g34980);
  dff DFF_1425(CK,RST,g2907,g34617);
  dff DFF_1426(CK,RST,g2912,g34618);
  dff DFF_1427(CK,RST,g2922,g34619);
  dff DFF_1428(CK,RST,g2936,g34620);
  dff DFF_1429(CK,RST,g2950,g34621);
  dff DFF_1430(CK,RST,g2960,g34622);
  dff DFF_1431(CK,RST,g2970,g34623);
  dff DFF_1432(CK,RST,g2902,g34801);
  dff DFF_1433(CK,RST,g2917,g34802);
  dff DFF_1434(CK,RST,g2927,g34803);
  dff DFF_1435(CK,RST,g2941,g34806);
  dff DFF_1436(CK,RST,g2955,g34807);
  dff DFF_1437(CK,RST,g2965,g34808);
  dff DFF_1438(CK,RST,g2975,g34804);
  dff DFF_1439(CK,RST,g3003,g21726);
  dff DFF_1440(CK,RST,g5,g12833);
  dff DFF_1441(CK,RST,g6,g34589);
  dff DFF_1442(CK,RST,g7,g34590);
  dff DFF_1443(CK,RST,g8,g34591);
  dff DFF_1444(CK,RST,g9,g34592);
  dff DFF_1445(CK,RST,g16,g34593);
  dff DFF_1446(CK,RST,g19,g34594);
  dff DFF_1447(CK,RST,g28,g34595);
  dff DFF_1448(CK,RST,g31,g34596);
  dff DFF_1449(CK,RST,g34,g34877);
  dff DFF_1450(CK,RST,g12,g30326);
  dff DFF_1451(CK,RST,g22,g29209);
  dff DFF_1452(CK,RST,g25,g15048);
  not NOT_1453(I11617,g1);
  not NOT_1454(g6754,I11617);
  not NOT_1455(I11620,g1);
  not NOT_1456(g6755,I11620);
  not NOT_1457(I11623,g28);
  not NOT_1458(g6756,I11623);
  not NOT_1459(I11626,g31);
  not NOT_1460(g6767,I11626);
  not NOT_1461(I11629,g19);
  not NOT_1462(g6772,I11629);
  not NOT_1463(I11632,g16);
  not NOT_1464(g6782,I11632);
  not NOT_1465(I11635,g9);
  not NOT_1466(g6789,I11635);
  not NOT_1467(g6799,g199);
  not NOT_1468(g6800,g203);
  not NOT_1469(g6801,g391);
  not NOT_1470(g6802,g468);
  not NOT_1471(g6803,g496);
  not NOT_1472(g6804,g490);
  not NOT_1473(g6808,g554);
  not NOT_1474(g6809,g341);
  not NOT_1475(g6810,g723);
  not NOT_1476(g6811,g714);
  not NOT_1477(g6814,g632);
  not NOT_1478(g6815,g929);
  not NOT_1479(g6816,g933);
  not NOT_1480(g6817,g956);
  not NOT_1481(g6818,g976);
  not NOT_1482(g6819,g1046);
  not NOT_1483(g6820,g1070);
  not NOT_1484(I11655,g1246);
  not NOT_1485(g6821,I11655);
  not NOT_1486(g6825,g979);
  not NOT_1487(g6826,g218);
  not NOT_1488(g6827,g1277);
  not NOT_1489(g6828,g1300);
  not NOT_1490(g6829,g1319);
  not NOT_1491(g6830,g1389);
  not NOT_1492(g6831,g1413);
  not NOT_1493(I11665,g1589);
  not NOT_1494(g6832,I11665);
  not NOT_1495(g6836,g1322);
  not NOT_1496(g6837,g968);
  not NOT_1497(g6838,g1724);
  not NOT_1498(g6839,g1858);
  not NOT_1499(g6840,g1992);
  not NOT_1500(g6841,g2145);
  not NOT_1501(g6845,g2126);
  not NOT_1502(g6846,g2152);
  not NOT_1503(g6847,g2283);
  not NOT_1504(g6848,g2417);
  not NOT_1505(g6849,g2551);
  not NOT_1506(g6850,g2704);
  not NOT_1507(g6854,g2685);
  not NOT_1508(g6855,g2711);
  not NOT_1509(I11682,g2756);
  not NOT_1510(g6856,I11682);
  not NOT_1511(I11685,g117);
  not NOT_1512(g6867,I11685);
  not NOT_1513(I11688,g70);
  not NOT_1514(g6868,I11688);
  not NOT_1515(I11691,g36);
  not NOT_1516(g6869,I11691);
  not NOT_1517(g6870,g3089);
  not NOT_1518(g6873,g3151);
  not NOT_1519(g6874,g3143);
  not NOT_1520(I11697,g3352);
  not NOT_1521(g6875,I11697);
  not NOT_1522(g6887,g3333);
  not NOT_1523(I11701,g4164);
  not NOT_1524(g6888,I11701);
  not NOT_1525(g6895,g3288);
  not NOT_1526(g6900,g3440);
  not NOT_1527(g6903,g3502);
  not NOT_1528(g6904,g3494);
  not NOT_1529(I11708,g3703);
  not NOT_1530(g6905,I11708);
  not NOT_1531(g6917,g3684);
  not NOT_1532(g6918,g3639);
  not NOT_1533(g6923,g3791);
  not NOT_1534(g6926,g3853);
  not NOT_1535(g6927,g3845);
  not NOT_1536(I11716,g4054);
  not NOT_1537(g6928,I11716);
  not NOT_1538(g6940,g4035);
  not NOT_1539(g6941,g3990);
  not NOT_1540(I11721,g4145);
  not NOT_1541(g6946,I11721);
  not NOT_1542(g6953,g4157);
  not NOT_1543(g6954,g4138);
  not NOT_1544(I11726,g4273);
  not NOT_1545(g6955,I11726);
  not NOT_1546(g6956,g4242);
  not NOT_1547(g6957,g2932);
  not NOT_1548(g6958,g4372);
  not NOT_1549(g6959,g4420);
  not NOT_1550(g6960,g1);
  not NOT_1551(I11734,g4473);
  not NOT_1552(g6961,I11734);
  not NOT_1553(I11737,g4467);
  not NOT_1554(g6971,I11737);
  not NOT_1555(I11740,g4519);
  not NOT_1556(g6972,I11740);
  not NOT_1557(I11743,g4564);
  not NOT_1558(g6973,I11743);
  not NOT_1559(I11746,g4570);
  not NOT_1560(g6974,I11746);
  not NOT_1561(g6975,g4507);
  not NOT_1562(I11750,g4474);
  not NOT_1563(g6976,I11750);
  not NOT_1564(I11753,g4492);
  not NOT_1565(g6977,I11753);
  not NOT_1566(g6978,g4616);
  not NOT_1567(g6982,g4531);
  not NOT_1568(g6983,g4698);
  not NOT_1569(g6984,g4709);
  not NOT_1570(g6985,g4669);
  not NOT_1571(g6986,g4743);
  not NOT_1572(g6987,g4754);
  not NOT_1573(g6988,g4765);
  not NOT_1574(g6989,g4575);
  not NOT_1575(g6990,g4742);
  not NOT_1576(g6991,g4888);
  not NOT_1577(g6992,g4899);
  not NOT_1578(g6993,g4859);
  not NOT_1579(g6994,g4933);
  not NOT_1580(g6995,g4944);
  not NOT_1581(g6996,g4955);
  not NOT_1582(g6997,g4578);
  not NOT_1583(g6998,g4932);
  not NOT_1584(g6999,g86);
  not NOT_1585(g7002,g5160);
  not NOT_1586(g7003,g5152);
  not NOT_1587(I11777,g5357);
  not NOT_1588(g7004,I11777);
  not NOT_1589(g7017,g128);
  not NOT_1590(g7018,g5297);
  not NOT_1591(g7023,g5445);
  not NOT_1592(g7026,g5507);
  not NOT_1593(g7027,g5499);
  not NOT_1594(I11785,g5703);
  not NOT_1595(g7028,I11785);
  not NOT_1596(g7040,g4821);
  not NOT_1597(g7041,g5644);
  not NOT_1598(g7046,g5791);
  not NOT_1599(g7049,g5853);
  not NOT_1600(g7050,g5845);
  not NOT_1601(I11793,g6049);
  not NOT_1602(g7051,I11793);
  not NOT_1603(g7063,g4831);
  not NOT_1604(g7064,g5990);
  not NOT_1605(g7069,g6137);
  not NOT_1606(g7072,g6199);
  not NOT_1607(g7073,g6191);
  not NOT_1608(I11801,g6395);
  not NOT_1609(g7074,I11801);
  not NOT_1610(g7086,g4826);
  not NOT_1611(g7087,g6336);
  not NOT_1612(g7092,g6483);
  not NOT_1613(g7095,g6545);
  not NOT_1614(g7096,g6537);
  not NOT_1615(I11809,g6741);
  not NOT_1616(g7097,I11809);
  not NOT_1617(g7109,g5011);
  not NOT_1618(g7110,g6682);
  not NOT_1619(g7115,g12);
  not NOT_1620(g7116,g22);
  not NOT_1621(I11816,g93);
  not NOT_1622(g7117,I11816);
  not NOT_1623(g7118,g832);
  not NOT_1624(I11820,g3869);
  not NOT_1625(g7121,I11820);
  not NOT_1626(g7132,g4558);
  not NOT_1627(g7134,g5029);
  not NOT_1628(g7138,g5360);
  not NOT_1629(I11835,g101);
  not NOT_1630(g7148,I11835);
  not NOT_1631(g7149,g4564);
  not NOT_1632(g7153,g5373);
  not NOT_1633(g7157,g5706);
  not NOT_1634(I11843,g111);
  not NOT_1635(g7161,I11843);
  not NOT_1636(g7162,g4521);
  not NOT_1637(g7163,g4593);
  not NOT_1638(g7166,g4311);
  not NOT_1639(g7170,g5719);
  not NOT_1640(g7174,g6052);
  not NOT_1641(g7178,g4392);
  not NOT_1642(g7183,g4608);
  not NOT_1643(g7187,g6065);
  not NOT_1644(g7191,g6398);
  not NOT_1645(g7195,g25);
  not NOT_1646(I11860,g43);
  not NOT_1647(g7196,I11860);
  not NOT_1648(g7197,g812);
  not NOT_1649(g7202,g4639);
  not NOT_1650(g7212,g6411);
  not NOT_1651(g7216,g822);
  not NOT_1652(g7219,g4405);
  not NOT_1653(g7222,g4427);
  not NOT_1654(g7224,g4601);
  not NOT_1655(g7231,g5);
  not NOT_1656(g7232,g4411);
  not NOT_1657(g7235,g4521);
  not NOT_1658(g7236,g4608);
  not NOT_1659(g7239,g5033);
  not NOT_1660(I11892,g4408);
  not NOT_1661(g7243,I11892);
  not NOT_1662(g7244,g4408);
  not NOT_1663(I11896,g4446);
  not NOT_1664(g7245,I11896);
  not NOT_1665(g7246,g4446);
  not NOT_1666(g7247,g5377);
  not NOT_1667(g7252,g1592);
  not NOT_1668(I11903,g4414);
  not NOT_1669(g7257,I11903);
  not NOT_1670(g7258,g4414);
  not NOT_1671(g7259,g4375);
  not NOT_1672(I11908,g4449);
  not NOT_1673(g7260,I11908);
  not NOT_1674(g7261,g4449);
  not NOT_1675(g7262,g5723);
  not NOT_1676(g7266,g35);
  not NOT_1677(g7267,g1604);
  not NOT_1678(g7268,g1636);
  not NOT_1679(g7275,g1728);
  not NOT_1680(g7280,g2153);
  not NOT_1681(g7285,g4643);
  not NOT_1682(g7289,g4382);
  not NOT_1683(g7293,g4452);
  not NOT_1684(g7296,g5313);
  not NOT_1685(g7297,g6069);
  not NOT_1686(g7301,g925);
  not NOT_1687(g7308,g1668);
  not NOT_1688(g7314,g1740);
  not NOT_1689(g7315,g1772);
  not NOT_1690(g7322,g1862);
  not NOT_1691(g7327,g2165);
  not NOT_1692(g7328,g2197);
  not NOT_1693(g7335,g2287);
  not NOT_1694(g7340,g4443);
  not NOT_1695(g7343,g5290);
  not NOT_1696(g7344,g5659);
  not NOT_1697(g7345,g6415);
  not NOT_1698(g7349,g1270);
  not NOT_1699(g7356,g1802);
  not NOT_1700(g7361,g1874);
  not NOT_1701(g7362,g1906);
  not NOT_1702(g7369,g1996);
  not NOT_1703(g7374,g2227);
  not NOT_1704(g7379,g2299);
  not NOT_1705(g7380,g2331);
  not NOT_1706(g7387,g2421);
  not NOT_1707(g7392,g4438);
  not NOT_1708(g7393,g5320);
  not NOT_1709(g7394,g5637);
  not NOT_1710(g7395,g6005);
  not NOT_1711(g7397,g890);
  not NOT_1712(g7400,g911);
  not NOT_1713(g7405,g1936);
  not NOT_1714(g7410,g2008);
  not NOT_1715(g7411,g2040);
  not NOT_1716(g7418,g2361);
  not NOT_1717(g7423,g2433);
  not NOT_1718(g7424,g2465);
  not NOT_1719(g7431,g2555);
  not NOT_1720(g7436,g5276);
  not NOT_1721(g7437,g5666);
  not NOT_1722(g7438,g5983);
  not NOT_1723(g7439,g6351);
  not NOT_1724(g7440,g329);
  not NOT_1725(g7441,g862);
  not NOT_1726(g7443,g914);
  not NOT_1727(g7446,g1256);
  not NOT_1728(g7451,g2070);
  not NOT_1729(g7456,g2495);
  not NOT_1730(g7461,g2567);
  not NOT_1731(g7462,g2599);
  not NOT_1732(g7470,g5623);
  not NOT_1733(g7471,g6012);
  not NOT_1734(g7472,g6329);
  not NOT_1735(g7473,g6697);
  not NOT_1736(I11980,g66);
  not NOT_1737(g7474,I11980);
  not NOT_1738(g7475,g896);
  not NOT_1739(g7479,g1008);
  not NOT_1740(g7487,g1259);
  not NOT_1741(g7490,g2629);
  not NOT_1742(g7495,g4375);
  not NOT_1743(g7496,g5969);
  not NOT_1744(g7497,g6358);
  not NOT_1745(g7498,g6675);
  not NOT_1746(I11992,g763);
  not NOT_1747(g7502,I11992);
  not NOT_1748(g7503,g1351);
  not NOT_1749(g7512,g5283);
  not NOT_1750(g7513,g6315);
  not NOT_1751(g7514,g6704);
  not NOT_1752(I12000,g582);
  not NOT_1753(g7515,I12000);
  not NOT_1754(I12003,g767);
  not NOT_1755(g7516,I12003);
  not NOT_1756(g7517,g962);
  not NOT_1757(g7518,g1024);
  not NOT_1758(g7519,g1157);
  not NOT_1759(g7521,g5630);
  not NOT_1760(g7522,g6661);
  not NOT_1761(g7523,g305);
  not NOT_1762(I12013,g590);
  not NOT_1763(g7526,I12013);
  not NOT_1764(I12016,g772);
  not NOT_1765(g7527,I12016);
  not NOT_1766(g7528,g930);
  not NOT_1767(g7532,g1157);
  not NOT_1768(g7533,g1306);
  not NOT_1769(g7534,g1367);
  not NOT_1770(g7535,g1500);
  not NOT_1771(g7536,g5976);
  not NOT_1772(g7537,g311);
  not NOT_1773(I12026,g344);
  not NOT_1774(g7540,I12026);
  not NOT_1775(g7541,g344);
  not NOT_1776(I12030,g595);
  not NOT_1777(g7542,I12030);
  not NOT_1778(I12033,g776);
  not NOT_1779(g7543,I12033);
  not NOT_1780(g7544,g918);
  not NOT_1781(g7548,g1036);
  not NOT_1782(g7553,g1274);
  not NOT_1783(g7557,g1500);
  not NOT_1784(I12041,g2741);
  not NOT_1785(g7558,I12041);
  not NOT_1786(g7563,g6322);
  not NOT_1787(g7564,g336);
  not NOT_1788(I12046,g613);
  not NOT_1789(g7565,I12046);
  not NOT_1790(I12049,g781);
  not NOT_1791(g7566,I12049);
  not NOT_1792(g7577,g1263);
  not NOT_1793(g7581,g1379);
  not NOT_1794(I12056,g2748);
  not NOT_1795(g7586,I12056);
  not NOT_1796(g7591,g6668);
  not NOT_1797(g7592,g347);
  not NOT_1798(I12061,g562);
  not NOT_1799(g7593,I12061);
  not NOT_1800(I12064,g617);
  not NOT_1801(g7594,I12064);
  not NOT_1802(I12067,g739);
  not NOT_1803(g7595,I12067);
  not NOT_1804(I12070,g785);
  not NOT_1805(g7596,I12070);
  not NOT_1806(g7597,g952);
  not NOT_1807(I12083,g568);
  not NOT_1808(g7615,I12083);
  not NOT_1809(I12086,g622);
  not NOT_1810(g7616,I12086);
  not NOT_1811(I12089,g744);
  not NOT_1812(g7617,I12089);
  not NOT_1813(I12092,g790);
  not NOT_1814(g7618,I12092);
  not NOT_1815(g7619,g1296);
  not NOT_1816(I12103,g572);
  not NOT_1817(g7623,I12103);
  not NOT_1818(I12106,g626);
  not NOT_1819(g7624,I12106);
  not NOT_1820(I12109,g749);
  not NOT_1821(g7625,I12109);
  not NOT_1822(I12112,g794);
  not NOT_1823(g7626,I12112);
  not NOT_1824(g7627,g4311);
  not NOT_1825(g7631,g74);
  not NOT_1826(I12117,g586);
  not NOT_1827(g7632,I12117);
  not NOT_1828(I12120,g632);
  not NOT_1829(g7633,I12120);
  not NOT_1830(I12123,g758);
  not NOT_1831(g7634,I12123);
  not NOT_1832(g7635,g1002);
  not NOT_1833(g7636,g4098);
  not NOT_1834(I12128,g4253);
  not NOT_1835(g7640,I12128);
  not NOT_1836(g7643,g4322);
  not NOT_1837(I12132,g577);
  not NOT_1838(g7647,I12132);
  not NOT_1839(I12135,g807);
  not NOT_1840(g7648,I12135);
  not NOT_1841(g7649,g1345);
  not NOT_1842(g7650,g4064);
  not NOT_1843(g7655,g4332);
  not NOT_1844(I12141,g599);
  not NOT_1845(g7659,I12141);
  not NOT_1846(I12144,g554);
  not NOT_1847(g7660,I12144);
  not NOT_1848(g7666,g4076);
  not NOT_1849(g7670,g4104);
  not NOT_1850(I12151,g604);
  not NOT_1851(g7674,I12151);
  not NOT_1852(g7680,g4108);
  not NOT_1853(g7686,g4659);
  not NOT_1854(I12159,g608);
  not NOT_1855(g7689,I12159);
  not NOT_1856(g7693,g4849);
  not NOT_1857(g7697,g4087);
  not NOT_1858(I12167,g5176);
  not NOT_1859(g7704,I12167);
  not NOT_1860(g7715,g1178);
  not NOT_1861(g7716,g1199);
  not NOT_1862(I12172,g2715);
  not NOT_1863(g7717,I12172);
  not NOT_1864(g7733,g4093);
  not NOT_1865(I12176,g5523);
  not NOT_1866(g7738,I12176);
  not NOT_1867(g7749,g996);
  not NOT_1868(g7750,g1070);
  not NOT_1869(g7751,g1521);
  not NOT_1870(g7752,g1542);
  not NOT_1871(I12183,g2719);
  not NOT_1872(g7753,I12183);
  not NOT_1873(g7765,g4165);
  not NOT_1874(I12189,g5869);
  not NOT_1875(g7766,I12189);
  not NOT_1876(g7778,g1339);
  not NOT_1877(g7779,g1413);
  not NOT_1878(g7780,g2878);
  not NOT_1879(g7785,g4621);
  not NOT_1880(g7788,g4674);
  not NOT_1881(I12199,g6215);
  not NOT_1882(g7791,I12199);
  not NOT_1883(g7802,g324);
  not NOT_1884(g7805,g4366);
  not NOT_1885(g7806,g4681);
  not NOT_1886(g7809,g4864);
  not NOT_1887(I12214,g6561);
  not NOT_1888(g7812,I12214);
  not NOT_1889(g7824,g4169);
  not NOT_1890(g7827,g4688);
  not NOT_1891(g7828,g4871);
  not NOT_1892(I12227,g34);
  not NOT_1893(g7831,I12227);
  not NOT_1894(g7835,g4125);
  not NOT_1895(g7840,g4878);
  not NOT_1896(g7841,g904);
  not NOT_1897(g7845,g1146);
  not NOT_1898(g7851,g921);
  not NOT_1899(g7854,g1152);
  not NOT_1900(g7858,g947);
  not NOT_1901(g7863,g1249);
  not NOT_1902(g7867,g1489);
  not NOT_1903(g7868,g1099);
  not NOT_1904(g7870,g1193);
  not NOT_1905(g7873,g1266);
  not NOT_1906(g7876,g1495);
  not NOT_1907(g7880,g1291);
  not NOT_1908(g7886,g1442);
  not NOT_1909(g7888,g1536);
  not NOT_1910(g7891,g2994);
  not NOT_1911(g7892,g4801);
  not NOT_1912(g7898,g4991);
  not NOT_1913(g7903,g969);
  not NOT_1914(g7907,g3072);
  not NOT_1915(g7908,g4157);
  not NOT_1916(g7909,g936);
  not NOT_1917(g7913,g1052);
  not NOT_1918(I12300,g1157);
  not NOT_1919(g7916,I12300);
  not NOT_1920(g7917,g1157);
  not NOT_1921(g7922,g1312);
  not NOT_1922(g7926,g3423);
  not NOT_1923(g7927,g4064);
  not NOT_1924(g7928,g4776);
  not NOT_1925(g7933,g907);
  not NOT_1926(g7936,g1061);
  not NOT_1927(g7939,g1280);
  not NOT_1928(g7943,g1395);
  not NOT_1929(I12314,g1500);
  not NOT_1930(g7946,I12314);
  not NOT_1931(g7947,g1500);
  not NOT_1932(g7952,g3774);
  not NOT_1933(g7953,g4966);
  not NOT_1934(g7957,g1252);
  not NOT_1935(g7960,g1404);
  not NOT_1936(g7963,g4146);
  not NOT_1937(g7964,g3155);
  not NOT_1938(g7970,g4688);
  not NOT_1939(g7971,g4818);
  not NOT_1940(g7972,g1046);
  not NOT_1941(g7975,g3040);
  not NOT_1942(g7980,g3161);
  not NOT_1943(g7985,g3506);
  not NOT_1944(g7991,g4878);
  not NOT_1945(g7992,g5008);
  not NOT_1946(I12333,g45);
  not NOT_1947(g7993,I12333);
  not NOT_1948(I12336,g52);
  not NOT_1949(g7994,I12336);
  not NOT_1950(g7995,g153);
  not NOT_1951(g7998,g392);
  not NOT_1952(g8002,g1389);
  not NOT_1953(g8005,g3025);
  not NOT_1954(g8009,g3106);
  not NOT_1955(g8011,g3167);
  not NOT_1956(g8016,g3391);
  not NOT_1957(g8021,g3512);
  not NOT_1958(g8026,g3857);
  not NOT_1959(I12355,g46);
  not NOT_1960(g8032,I12355);
  not NOT_1961(g8033,g157);
  not NOT_1962(g8037,g405);
  not NOT_1963(I12360,g528);
  not NOT_1964(g8038,I12360);
  not NOT_1965(g8046,g528);
  not NOT_1966(g8052,g1211);
  not NOT_1967(g8055,g1236);
  not NOT_1968(g8056,g1246);
  not NOT_1969(g8057,g3068);
  not NOT_1970(g8058,g3115);
  not NOT_1971(g8059,g3171);
  not NOT_1972(g8064,g3376);
  not NOT_1973(g8068,g3457);
  not NOT_1974(g8070,g3518);
  not NOT_1975(g8075,g3742);
  not NOT_1976(g8080,g3863);
  not NOT_1977(I12382,g47);
  not NOT_1978(g8085,I12382);
  not NOT_1979(g8087,g1157);
  not NOT_1980(g8088,g1554);
  not NOT_1981(g8091,g1579);
  not NOT_1982(g8092,g1589);
  not NOT_1983(g8093,g1624);
  not NOT_1984(g8097,g3029);
  not NOT_1985(g8102,g3072);
  not NOT_1986(g8106,g3133);
  not NOT_1987(g8107,g3179);
  not NOT_1988(g8112,g3419);
  not NOT_1989(g8113,g3466);
  not NOT_1990(g8114,g3522);
  not NOT_1991(g8119,g3727);
  not NOT_1992(g8123,g3808);
  not NOT_1993(g8125,g3869);
  not NOT_1994(g8130,g4515);
  not NOT_1995(I12411,g4809);
  not NOT_1996(g8132,I12411);
  not NOT_1997(g8133,g4809);
  not NOT_1998(I12415,g48);
  not NOT_1999(g8134,I12415);
  not NOT_2000(I12418,g55);
  not NOT_2001(g8135,I12418);
  not NOT_2002(g8136,g269);
  not NOT_2003(g8137,g411);
  not NOT_2004(g8138,g1500);
  not NOT_2005(g8139,g1648);
  not NOT_2006(g8146,g1760);
  not NOT_2007(g8150,g2185);
  not NOT_2008(g8154,g3139);
  not NOT_2009(g8155,g3380);
  not NOT_2010(g8160,g3423);
  not NOT_2011(g8164,g3484);
  not NOT_2012(g8165,g3530);
  not NOT_2013(g8170,g3770);
  not NOT_2014(g8171,g3817);
  not NOT_2015(g8172,g3873);
  not NOT_2016(I12437,g4999);
  not NOT_2017(g8178,I12437);
  not NOT_2018(g8179,g4999);
  not NOT_2019(g8180,g262);
  not NOT_2020(g8181,g424);
  not NOT_2021(g8183,g482);
  not NOT_2022(g8186,g990);
  not NOT_2023(g8187,g1657);
  not NOT_2024(g8195,g1783);
  not NOT_2025(g8201,g1894);
  not NOT_2026(g8205,g2208);
  not NOT_2027(g8211,g2319);
  not NOT_2028(I12451,g3092);
  not NOT_2029(g8215,I12451);
  not NOT_2030(g8216,g3092);
  not NOT_2031(g8217,g3143);
  not NOT_2032(g8218,g3490);
  not NOT_2033(g8219,g3731);
  not NOT_2034(g8224,g3774);
  not NOT_2035(g8228,g3835);
  not NOT_2036(g8229,g3881);
  not NOT_2037(I12463,g4812);
  not NOT_2038(g8235,I12463);
  not NOT_2039(g8236,g4812);
  not NOT_2040(g8237,g255);
  not NOT_2041(g8239,g1056);
  not NOT_2042(g8240,g1333);
  not NOT_2043(g8241,g1792);
  not NOT_2044(g8249,g1917);
  not NOT_2045(g8255,g2028);
  not NOT_2046(g8259,g2217);
  not NOT_2047(g8267,g2342);
  not NOT_2048(g8273,g2453);
  not NOT_2049(I12483,g3096);
  not NOT_2050(g8277,I12483);
  not NOT_2051(g8278,g3096);
  not NOT_2052(I12487,g3443);
  not NOT_2053(g8279,I12487);
  not NOT_2054(g8280,g3443);
  not NOT_2055(g8281,g3494);
  not NOT_2056(g8282,g3841);
  not NOT_2057(I12493,g5002);
  not NOT_2058(g8283,I12493);
  not NOT_2059(g8284,g5002);
  not NOT_2060(I12497,g49);
  not NOT_2061(g8285,I12497);
  not NOT_2062(g8286,g53);
  not NOT_2063(g8287,g160);
  not NOT_2064(g8290,g218);
  not NOT_2065(I12503,g215);
  not NOT_2066(g8291,I12503);
  not NOT_2067(g8296,g246);
  not NOT_2068(g8297,g142);
  not NOT_2069(g8300,g1242);
  not NOT_2070(g8301,g1399);
  not NOT_2071(g8302,g1926);
  not NOT_2072(g8310,g2051);
  not NOT_2073(g8316,g2351);
  not NOT_2074(g8324,g2476);
  not NOT_2075(g8330,g2587);
  not NOT_2076(g8334,g3034);
  not NOT_2077(g8340,g3050);
  not NOT_2078(g8341,g3119);
  not NOT_2079(I12519,g3447);
  not NOT_2080(g8342,I12519);
  not NOT_2081(g8343,g3447);
  not NOT_2082(I12523,g3794);
  not NOT_2083(g8344,I12523);
  not NOT_2084(g8345,g3794);
  not NOT_2085(g8346,g3845);
  not NOT_2086(g8350,g4646);
  not NOT_2087(I12530,g4815);
  not NOT_2088(g8353,I12530);
  not NOT_2089(g8354,g4815);
  not NOT_2090(I12534,g50);
  not NOT_2091(g8355,I12534);
  not NOT_2092(g8356,g54);
  not NOT_2093(I12538,g58);
  not NOT_2094(g8357,I12538);
  not NOT_2095(I12541,g194);
  not NOT_2096(g8358,I12541);
  not NOT_2097(g8362,g194);
  not NOT_2098(g8363,g239);
  not NOT_2099(g8364,g1585);
  not NOT_2100(g8365,g2060);
  not NOT_2101(g8373,g2485);
  not NOT_2102(g8381,g2610);
  not NOT_2103(g8387,g3080);
  not NOT_2104(g8388,g3010);
  not NOT_2105(g8389,g3125);
  not NOT_2106(g8390,g3385);
  not NOT_2107(g8396,g3401);
  not NOT_2108(g8397,g3470);
  not NOT_2109(I12563,g3798);
  not NOT_2110(g8398,I12563);
  not NOT_2111(g8399,g3798);
  not NOT_2112(g8400,g4836);
  not NOT_2113(I12568,g5005);
  not NOT_2114(g8403,I12568);
  not NOT_2115(g8404,g5005);
  not NOT_2116(I12572,g51);
  not NOT_2117(g8405,I12572);
  not NOT_2118(g8406,g232);
  not NOT_2119(g8407,g1171);
  not NOT_2120(I12577,g1227);
  not NOT_2121(g8411,I12577);
  not NOT_2122(I12580,g1239);
  not NOT_2123(g8416,I12580);
  not NOT_2124(g8418,g2619);
  not NOT_2125(g8426,g3045);
  not NOT_2126(g8431,g3085);
  not NOT_2127(g8438,g3100);
  not NOT_2128(g8439,g3129);
  not NOT_2129(g8440,g3431);
  not NOT_2130(g8441,g3361);
  not NOT_2131(g8442,g3476);
  not NOT_2132(g8443,g3736);
  not NOT_2133(g8449,g3752);
  not NOT_2134(g8450,g3821);
  not NOT_2135(g8451,g4057);
  not NOT_2136(g8456,g56);
  not NOT_2137(g8457,g225);
  not NOT_2138(g8458,g294);
  not NOT_2139(g8462,g1183);
  not NOT_2140(g8466,g1514);
  not NOT_2141(I12605,g1570);
  not NOT_2142(g8470,I12605);
  not NOT_2143(I12608,g1582);
  not NOT_2144(g8475,I12608);
  not NOT_2145(g8477,g3061);
  not NOT_2146(g8478,g3103);
  not NOT_2147(g8479,g3057);
  not NOT_2148(g8480,g3147);
  not NOT_2149(I12618,g3338);
  not NOT_2150(g8481,I12618);
  not NOT_2151(g8492,g3396);
  not NOT_2152(g8497,g3436);
  not NOT_2153(g8504,g3451);
  not NOT_2154(g8505,g3480);
  not NOT_2155(g8506,g3782);
  not NOT_2156(g8507,g3712);
  not NOT_2157(g8508,g3827);
  not NOT_2158(g8509,g4141);
  not NOT_2159(g8514,g4258);
  not NOT_2160(I12631,g1242);
  not NOT_2161(g8515,I12631);
  not NOT_2162(g8519,g287);
  not NOT_2163(g8522,g298);
  not NOT_2164(g8526,g1526);
  not NOT_2165(g8531,g3288);
  not NOT_2166(g8534,g3338);
  not NOT_2167(g8538,g3412);
  not NOT_2168(g8539,g3454);
  not NOT_2169(g8540,g3408);
  not NOT_2170(g8541,g3498);
  not NOT_2171(I12644,g3689);
  not NOT_2172(g8542,I12644);
  not NOT_2173(g8553,g3747);
  not NOT_2174(g8558,g3787);
  not NOT_2175(g8565,g3802);
  not NOT_2176(g8566,g3831);
  not NOT_2177(g8567,g4082);
  not NOT_2178(g8571,g57);
  not NOT_2179(I12654,g1585);
  not NOT_2180(g8572,I12654);
  not NOT_2181(g8575,g291);
  not NOT_2182(g8579,g2771);
  not NOT_2183(g8584,g3639);
  not NOT_2184(g8587,g3689);
  not NOT_2185(g8591,g3763);
  not NOT_2186(g8592,g3805);
  not NOT_2187(g8593,g3759);
  not NOT_2188(g8594,g3849);
  not NOT_2189(I12666,g4040);
  not NOT_2190(g8595,I12666);
  not NOT_2191(g8606,g4653);
  not NOT_2192(g8607,g37);
  not NOT_2193(g8608,g278);
  not NOT_2194(g8612,g2775);
  not NOT_2195(g8616,g2803);
  not NOT_2196(g8620,g3065);
  not NOT_2197(g8623,g3990);
  not NOT_2198(g8626,g4040);
  not NOT_2199(g8630,g4843);
  not NOT_2200(g8631,g283);
  not NOT_2201(g8635,g2783);
  not NOT_2202(g8639,g2807);
  not NOT_2203(g8644,g3352);
  not NOT_2204(g8647,g3416);
  not NOT_2205(g8650,g4664);
  not NOT_2206(g8651,g758);
  not NOT_2207(g8654,g1087);
  not NOT_2208(g8655,g2787);
  not NOT_2209(g8659,g2815);
  not NOT_2210(g8663,g3343);
  not NOT_2211(g8666,g3703);
  not NOT_2212(g8669,g3767);
  not NOT_2213(g8672,g4669);
  not NOT_2214(g8673,g4737);
  not NOT_2215(g8676,g4821);
  not NOT_2216(g8677,g4854);
  not NOT_2217(g8680,g686);
  not NOT_2218(g8681,g763);
  not NOT_2219(g8685,g1430);
  not NOT_2220(g8686,g2819);
  not NOT_2221(g8696,g3347);
  not NOT_2222(g8697,g3694);
  not NOT_2223(g8700,g4054);
  not NOT_2224(I12709,g4284);
  not NOT_2225(g8703,I12709);
  not NOT_2226(I12712,g59);
  not NOT_2227(g8712,I12712);
  not NOT_2228(g8713,g4826);
  not NOT_2229(g8714,g4859);
  not NOT_2230(g8715,g4927);
  not NOT_2231(g8718,g3333);
  not NOT_2232(I12719,g365);
  not NOT_2233(g8719,I12719);
  not NOT_2234(g8725,g739);
  not NOT_2235(g8733,g3698);
  not NOT_2236(g8734,g4045);
  not NOT_2237(I12735,g4572);
  not NOT_2238(g8740,I12735);
  not NOT_2239(g8741,g4821);
  not NOT_2240(g8742,g4035);
  not NOT_2241(g8743,g550);
  not NOT_2242(g8744,g691);
  not NOT_2243(g8745,g744);
  not NOT_2244(g8748,g776);
  not NOT_2245(g8756,g4049);
  not NOT_2246(I12746,g4087);
  not NOT_2247(g8757,I12746);
  not NOT_2248(I12749,g4575);
  not NOT_2249(g8763,I12749);
  not NOT_2250(g8764,g4826);
  not NOT_2251(g8765,g3333);
  not NOT_2252(g8766,g572);
  not NOT_2253(g8770,g749);
  not NOT_2254(g8774,g781);
  not NOT_2255(I12758,g4093);
  not NOT_2256(g8778,I12758);
  not NOT_2257(I12761,g4188);
  not NOT_2258(g8783,I12761);
  not NOT_2259(I12764,g4194);
  not NOT_2260(g8784,I12764);
  not NOT_2261(I12767,g4197);
  not NOT_2262(g8785,I12767);
  not NOT_2263(I12770,g4200);
  not NOT_2264(g8786,I12770);
  not NOT_2265(I12773,g4204);
  not NOT_2266(g8787,I12773);
  not NOT_2267(I12776,g4207);
  not NOT_2268(g8788,I12776);
  not NOT_2269(I12779,g4210);
  not NOT_2270(g8789,I12779);
  not NOT_2271(I12787,g4311);
  not NOT_2272(g8791,I12787);
  not NOT_2273(I12790,g4340);
  not NOT_2274(g8792,I12790);
  not NOT_2275(I12793,g4578);
  not NOT_2276(g8795,I12793);
  not NOT_2277(g8796,g4785);
  not NOT_2278(g8804,g4035);
  not NOT_2279(I12799,g59);
  not NOT_2280(g8805,I12799);
  not NOT_2281(g8807,g79);
  not NOT_2282(g8808,g595);
  not NOT_2283(I12805,g4098);
  not NOT_2284(g8812,I12805);
  not NOT_2285(I12808,g4322);
  not NOT_2286(g8818,I12808);
  not NOT_2287(I12811,g4340);
  not NOT_2288(g8821,I12811);
  not NOT_2289(g8822,g4975);
  not NOT_2290(g8830,g767);
  not NOT_2291(g8833,g794);
  not NOT_2292(g8836,g736);
  not NOT_2293(I12819,g4277);
  not NOT_2294(g8839,I12819);
  not NOT_2295(g8840,g4277);
  not NOT_2296(I12823,g4311);
  not NOT_2297(g8841,I12823);
  not NOT_2298(I12826,g4349);
  not NOT_2299(g8844,I12826);
  not NOT_2300(g8848,g358);
  not NOT_2301(g8851,g590);
  not NOT_2302(g8854,g613);
  not NOT_2303(g8858,g671);
  not NOT_2304(g8859,g772);
  not NOT_2305(I12837,g4222);
  not NOT_2306(g8870,I12837);
  not NOT_2307(g8872,g4258);
  not NOT_2308(I12855,g4311);
  not NOT_2309(g8876,I12855);
  not NOT_2310(I12858,g4340);
  not NOT_2311(g8879,I12858);
  not NOT_2312(I12861,g4372);
  not NOT_2313(g8880,I12861);
  not NOT_2314(g8883,g4709);
  not NOT_2315(g8890,g376);
  not NOT_2316(g8891,g582);
  not NOT_2317(g8895,g599);
  not NOT_2318(g8898,g676);
  not NOT_2319(g8899,g807);
  not NOT_2320(g8903,g1075);
  not NOT_2321(g8912,g4180);
  not NOT_2322(g8914,g4264);
  not NOT_2323(I12884,g4213);
  not NOT_2324(g8915,I12884);
  not NOT_2325(I12887,g4216);
  not NOT_2326(g8916,I12887);
  not NOT_2327(I12890,g4219);
  not NOT_2328(g8917,I12890);
  not NOT_2329(I12893,g4226);
  not NOT_2330(g8918,I12893);
  not NOT_2331(I12896,g4229);
  not NOT_2332(g8919,I12896);
  not NOT_2333(I12899,g4232);
  not NOT_2334(g8920,I12899);
  not NOT_2335(I12907,g4322);
  not NOT_2336(g8922,I12907);
  not NOT_2337(I12910,g4340);
  not NOT_2338(g8925,I12910);
  not NOT_2339(g8928,g4340);
  not NOT_2340(g8938,g4899);
  not NOT_2341(g8944,g370);
  not NOT_2342(g8945,g608);
  not NOT_2343(g8948,g785);
  not NOT_2344(g8951,g554);
  not NOT_2345(g8954,g1079);
  not NOT_2346(g8955,g1418);
  not NOT_2347(g8964,g4269);
  not NOT_2348(I12927,g4332);
  not NOT_2349(g8971,I12927);
  not NOT_2350(I12930,g4349);
  not NOT_2351(g8974,I12930);
  not NOT_2352(g8977,g4349);
  not NOT_2353(I12935,g6753);
  not NOT_2354(g8989,I12935);
  not NOT_2355(g8990,g146);
  not NOT_2356(g8993,g385);
  not NOT_2357(g8997,g577);
  not NOT_2358(g9000,g632);
  not NOT_2359(g9003,g790);
  not NOT_2360(g9007,g1083);
  not NOT_2361(g9011,g1422);
  not NOT_2362(g9014,g3004);
  not NOT_2363(g9018,g4273);
  not NOT_2364(I12950,g4287);
  not NOT_2365(g9019,I12950);
  not NOT_2366(g9020,g4287);
  not NOT_2367(I12954,g4358);
  not NOT_2368(g9021,I12954);
  not NOT_2369(g9024,g4358);
  not NOT_2370(g9030,g4793);
  not NOT_2371(g9036,g5084);
  not NOT_2372(g9037,g164);
  not NOT_2373(g9040,g499);
  not NOT_2374(g9044,g604);
  not NOT_2375(I12963,g640);
  not NOT_2376(g9048,I12963);
  not NOT_2377(g9049,g640);
  not NOT_2378(g9050,g1087);
  not NOT_2379(g9051,g1426);
  not NOT_2380(g9056,g3017);
  not NOT_2381(g9060,g3355);
  not NOT_2382(g9064,g4983);
  not NOT_2383(g9070,g5428);
  not NOT_2384(g9071,g2831);
  not NOT_2385(g9072,g2994);
  not NOT_2386(g9073,g150);
  not NOT_2387(g9077,g504);
  not NOT_2388(g9083,g626);
  not NOT_2389(g9086,g847);
  not NOT_2390(g9091,g1430);
  not NOT_2391(g9095,g3368);
  not NOT_2392(g9099,g3706);
  not NOT_2393(g9103,g5774);
  not NOT_2394(I12987,g12);
  not NOT_2395(g9104,I12987);
  not NOT_2396(g9152,g2834);
  not NOT_2397(I12991,g6752);
  not NOT_2398(g9153,I12991);
  not NOT_2399(I12994,g6748);
  not NOT_2400(g9154,I12994);
  not NOT_2401(I12997,g351);
  not NOT_2402(g9155,I12997);
  not NOT_2403(g9158,g513);
  not NOT_2404(g9162,g622);
  not NOT_2405(g9166,g837);
  not NOT_2406(g9174,g1205);
  not NOT_2407(g9180,g3719);
  not NOT_2408(g9184,g6120);
  not NOT_2409(I13007,g65);
  not NOT_2410(g9185,I13007);
  not NOT_2411(I13010,g6749);
  not NOT_2412(g9186,I13010);
  not NOT_2413(g9187,g518);
  not NOT_2414(g9194,g827);
  not NOT_2415(g9197,g1221);
  not NOT_2416(g9200,g1548);
  not NOT_2417(g9206,g5164);
  not NOT_2418(g9212,g6466);
  not NOT_2419(I13020,g6750);
  not NOT_2420(g9213,I13020);
  not NOT_2421(g9214,g617);
  not NOT_2422(g9220,g843);
  not NOT_2423(g9223,g1216);
  not NOT_2424(g9226,g1564);
  not NOT_2425(g9229,g5052);
  not NOT_2426(g9234,g5170);
  not NOT_2427(g9239,g5511);
  not NOT_2428(I13031,g6747);
  not NOT_2429(g9245,I13031);
  not NOT_2430(g9247,g1559);
  not NOT_2431(g9250,g1600);
  not NOT_2432(I13037,g4304);
  not NOT_2433(g9251,I13037);
  not NOT_2434(g9252,g4304);
  not NOT_2435(g9253,g5037);
  not NOT_2436(g9257,g5115);
  not NOT_2437(g9259,g5176);
  not NOT_2438(g9264,g5396);
  not NOT_2439(g9269,g5517);
  not NOT_2440(g9274,g5857);
  not NOT_2441(I13054,g6744);
  not NOT_2442(g9280,I13054);
  not NOT_2443(I13057,g112);
  not NOT_2444(g9281,I13057);
  not NOT_2445(g9282,g723);
  not NOT_2446(g9283,g1736);
  not NOT_2447(g9284,g2161);
  not NOT_2448(g9285,g2715);
  not NOT_2449(g9291,g3021);
  not NOT_2450(g9298,g5080);
  not NOT_2451(g9299,g5124);
  not NOT_2452(g9300,g5180);
  not NOT_2453(g9305,g5381);
  not NOT_2454(g9309,g5462);
  not NOT_2455(g9311,g5523);
  not NOT_2456(g9316,g5742);
  not NOT_2457(g9321,g5863);
  not NOT_2458(g9326,g6203);
  not NOT_2459(g9332,g64);
  not NOT_2460(g9333,g417);
  not NOT_2461(g9337,g1608);
  not NOT_2462(g9338,g1870);
  not NOT_2463(g9339,g2295);
  not NOT_2464(I13094,g2724);
  not NOT_2465(g9340,I13094);
  not NOT_2466(g9354,g2719);
  not NOT_2467(g9360,g3372);
  not NOT_2468(g9364,g5041);
  not NOT_2469(g9369,g5084);
  not NOT_2470(g9373,g5142);
  not NOT_2471(g9374,g5188);
  not NOT_2472(g9379,g5424);
  not NOT_2473(g9380,g5471);
  not NOT_2474(g9381,g5527);
  not NOT_2475(g9386,g5727);
  not NOT_2476(g9390,g5808);
  not NOT_2477(g9392,g5869);
  not NOT_2478(g9397,g6088);
  not NOT_2479(g9402,g6209);
  not NOT_2480(g9407,g6549);
  not NOT_2481(g9413,g1744);
  not NOT_2482(g9414,g2004);
  not NOT_2483(g9415,g2169);
  not NOT_2484(g9416,g2429);
  not NOT_2485(I13124,g2729);
  not NOT_2486(g9417,I13124);
  not NOT_2487(g9429,g3723);
  not NOT_2488(g9433,g5148);
  not NOT_2489(g9434,g5385);
  not NOT_2490(g9439,g5428);
  not NOT_2491(g9443,g5489);
  not NOT_2492(g9444,g5535);
  not NOT_2493(g9449,g5770);
  not NOT_2494(g9450,g5817);
  not NOT_2495(g9451,g5873);
  not NOT_2496(g9456,g6073);
  not NOT_2497(g9460,g6154);
  not NOT_2498(g9462,g6215);
  not NOT_2499(g9467,g6434);
  not NOT_2500(g9472,g6555);
  not NOT_2501(I13149,g6745);
  not NOT_2502(g9477,I13149);
  not NOT_2503(I13152,g6746);
  not NOT_2504(g9478,I13152);
  not NOT_2505(g9480,g559);
  not NOT_2506(g9484,g1612);
  not NOT_2507(g9488,g1878);
  not NOT_2508(g9489,g2303);
  not NOT_2509(g9490,g2563);
  not NOT_2510(g9491,g2729);
  not NOT_2511(g9492,g2759);
  not NOT_2512(g9496,g3303);
  not NOT_2513(I13166,g5101);
  not NOT_2514(g9497,I13166);
  not NOT_2515(g9498,g5101);
  not NOT_2516(g9499,g5152);
  not NOT_2517(g9500,g5495);
  not NOT_2518(g9501,g5731);
  not NOT_2519(g9506,g5774);
  not NOT_2520(g9510,g5835);
  not NOT_2521(g9511,g5881);
  not NOT_2522(g9516,g6116);
  not NOT_2523(g9517,g6163);
  not NOT_2524(g9518,g6219);
  not NOT_2525(g9523,g6419);
  not NOT_2526(g9527,g6500);
  not NOT_2527(g9529,g6561);
  not NOT_2528(g9534,g90);
  not NOT_2529(g9537,g1748);
  not NOT_2530(g9541,g2012);
  not NOT_2531(g9542,g2173);
  not NOT_2532(g9546,g2437);
  not NOT_2533(g9547,g2735);
  not NOT_2534(g9551,g3281);
  not NOT_2535(g9552,g3654);
  not NOT_2536(I13202,g5105);
  not NOT_2537(g9553,I13202);
  not NOT_2538(g9554,g5105);
  not NOT_2539(I13206,g5448);
  not NOT_2540(g9555,I13206);
  not NOT_2541(g9556,g5448);
  not NOT_2542(g9557,g5499);
  not NOT_2543(g9558,g5841);
  not NOT_2544(g9559,g6077);
  not NOT_2545(g9564,g6120);
  not NOT_2546(g9568,g6181);
  not NOT_2547(g9569,g6227);
  not NOT_2548(g9574,g6462);
  not NOT_2549(g9575,g6509);
  not NOT_2550(g9576,g6565);
  not NOT_2551(g9581,g91);
  not NOT_2552(g9582,g703);
  not NOT_2553(g9585,g1616);
  not NOT_2554(g9590,g1882);
  not NOT_2555(g9594,g2307);
  not NOT_2556(g9598,g2571);
  not NOT_2557(g9599,g3310);
  not NOT_2558(g9600,g3632);
  not NOT_2559(g9601,g4005);
  not NOT_2560(g9607,g5046);
  not NOT_2561(g9613,g5062);
  not NOT_2562(g9614,g5128);
  not NOT_2563(I13236,g5452);
  not NOT_2564(g9615,I13236);
  not NOT_2565(g9616,g5452);
  not NOT_2566(I13240,g5794);
  not NOT_2567(g9617,I13240);
  not NOT_2568(g9618,g5794);
  not NOT_2569(g9619,g5845);
  not NOT_2570(g9620,g6187);
  not NOT_2571(g9621,g6423);
  not NOT_2572(g9626,g6466);
  not NOT_2573(g9630,g6527);
  not NOT_2574(g9631,g6573);
  not NOT_2575(g9636,g72);
  not NOT_2576(I13252,g6751);
  not NOT_2577(g9637,I13252);
  not NOT_2578(g9638,g1620);
  not NOT_2579(g9639,g1752);
  not NOT_2580(g9644,g2016);
  not NOT_2581(g9648,g2177);
  not NOT_2582(g9653,g2441);
  not NOT_2583(g9657,g2763);
  not NOT_2584(g9660,g3267);
  not NOT_2585(g9661,g3661);
  not NOT_2586(g9662,g3983);
  not NOT_2587(g9669,g5092);
  not NOT_2588(g9670,g5022);
  not NOT_2589(g9671,g5134);
  not NOT_2590(g9672,g5390);
  not NOT_2591(g9678,g5406);
  not NOT_2592(g9679,g5475);
  not NOT_2593(I13276,g5798);
  not NOT_2594(g9680,I13276);
  not NOT_2595(g9681,g5798);
  not NOT_2596(I13280,g6140);
  not NOT_2597(g9682,I13280);
  not NOT_2598(g9683,g6140);
  not NOT_2599(g9684,g6191);
  not NOT_2600(g9685,g6533);
  not NOT_2601(g9686,g73);
  not NOT_2602(I13287,g110);
  not NOT_2603(g9687,I13287);
  not NOT_2604(g9688,g113);
  not NOT_2605(g9689,g124);
  not NOT_2606(g9690,g732);
  not NOT_2607(g9691,g1706);
  not NOT_2608(g9692,g1756);
  not NOT_2609(g9693,g1886);
  not NOT_2610(g9698,g2181);
  not NOT_2611(g9699,g2311);
  not NOT_2612(g9704,g2575);
  not NOT_2613(g9708,g2741);
  not NOT_2614(g9713,g3618);
  not NOT_2615(g9714,g4012);
  not NOT_2616(g9716,g5057);
  not NOT_2617(g9721,g5097);
  not NOT_2618(g9728,g5109);
  not NOT_2619(g9729,g5138);
  not NOT_2620(g9730,g5436);
  not NOT_2621(g9731,g5366);
  not NOT_2622(g9732,g5481);
  not NOT_2623(g9733,g5736);
  not NOT_2624(g9739,g5752);
  not NOT_2625(g9740,g5821);
  not NOT_2626(I13317,g6144);
  not NOT_2627(g9741,I13317);
  not NOT_2628(g9742,g6144);
  not NOT_2629(I13321,g6486);
  not NOT_2630(g9743,I13321);
  not NOT_2631(g9744,g6486);
  not NOT_2632(g9745,g6537);
  not NOT_2633(I13326,g66);
  not NOT_2634(g9746,I13326);
  not NOT_2635(I13329,g86);
  not NOT_2636(g9747,I13329);
  not NOT_2637(g9748,g114);
  not NOT_2638(g9749,g1691);
  not NOT_2639(g9751,g1710);
  not NOT_2640(g9752,g1840);
  not NOT_2641(g9753,g1890);
  not NOT_2642(g9754,g2020);
  not NOT_2643(g9759,g2265);
  not NOT_2644(g9760,g2315);
  not NOT_2645(g9761,g2445);
  not NOT_2646(g9766,g2748);
  not NOT_2647(g9771,g3969);
  not NOT_2648(I13352,g4146);
  not NOT_2649(g9772,I13352);
  not NOT_2650(g9776,g5073);
  not NOT_2651(g9777,g5112);
  not NOT_2652(g9778,g5069);
  not NOT_2653(g9779,g5156);
  not NOT_2654(I13360,g5343);
  not NOT_2655(g9780,I13360);
  not NOT_2656(g9792,g5401);
  not NOT_2657(g9797,g5441);
  not NOT_2658(g9804,g5456);
  not NOT_2659(g9805,g5485);
  not NOT_2660(g9806,g5782);
  not NOT_2661(g9807,g5712);
  not NOT_2662(g9808,g5827);
  not NOT_2663(g9809,g6082);
  not NOT_2664(g9815,g6098);
  not NOT_2665(g9816,g6167);
  not NOT_2666(I13374,g6490);
  not NOT_2667(g9817,I13374);
  not NOT_2668(g9818,g6490);
  not NOT_2669(g9819,g92);
  not NOT_2670(g9820,g99);
  not NOT_2671(g9821,g115);
  not NOT_2672(g9822,g125);
  not NOT_2673(g9824,g1825);
  not NOT_2674(g9826,g1844);
  not NOT_2675(g9827,g1974);
  not NOT_2676(g9828,g2024);
  not NOT_2677(g9829,g2250);
  not NOT_2678(g9831,g2269);
  not NOT_2679(g9832,g2399);
  not NOT_2680(g9833,g2449);
  not NOT_2681(g9834,g2579);
  not NOT_2682(g9839,g2724);
  not NOT_2683(g9842,g3274);
  not NOT_2684(g9843,g4311);
  not NOT_2685(g9848,g4462);
  not NOT_2686(g9853,g5297);
  not NOT_2687(g9856,g5343);
  not NOT_2688(g9860,g5417);
  not NOT_2689(g9861,g5459);
  not NOT_2690(g9862,g5413);
  not NOT_2691(g9863,g5503);
  not NOT_2692(I13424,g5689);
  not NOT_2693(g9864,I13424);
  not NOT_2694(g9875,g5747);
  not NOT_2695(g9880,g5787);
  not NOT_2696(g9887,g5802);
  not NOT_2697(g9888,g5831);
  not NOT_2698(g9889,g6128);
  not NOT_2699(g9890,g6058);
  not NOT_2700(g9891,g6173);
  not NOT_2701(g9892,g6428);
  not NOT_2702(g9898,g6444);
  not NOT_2703(g9899,g6513);
  not NOT_2704(g9900,g6);
  not NOT_2705(g9901,g84);
  not NOT_2706(g9902,g100);
  not NOT_2707(g9903,g681);
  not NOT_2708(g9905,g802);
  not NOT_2709(g9907,g1959);
  not NOT_2710(g9909,g1978);
  not NOT_2711(g9910,g2108);
  not NOT_2712(g9911,g2384);
  not NOT_2713(g9913,g2403);
  not NOT_2714(g9914,g2533);
  not NOT_2715(g9915,g2583);
  not NOT_2716(g9916,g3625);
  not NOT_2717(I13473,g4157);
  not NOT_2718(g9917,I13473);
  not NOT_2719(g9920,g4322);
  not NOT_2720(g9924,g5644);
  not NOT_2721(g9927,g5689);
  not NOT_2722(g9931,g5763);
  not NOT_2723(g9932,g5805);
  not NOT_2724(g9933,g5759);
  not NOT_2725(g9934,g5849);
  not NOT_2726(I13483,g6035);
  not NOT_2727(g9935,I13483);
  not NOT_2728(g9946,g6093);
  not NOT_2729(g9951,g6133);
  not NOT_2730(g9958,g6148);
  not NOT_2731(g9959,g6177);
  not NOT_2732(g9960,g6474);
  not NOT_2733(g9961,g6404);
  not NOT_2734(g9962,g6519);
  not NOT_2735(g9963,g7);
  not NOT_2736(g9964,g126);
  not NOT_2737(g9965,g127);
  not NOT_2738(g9969,g1682);
  not NOT_2739(g9970,g1714);
  not NOT_2740(g9971,g2093);
  not NOT_2741(g9973,g2112);
  not NOT_2742(g9974,g2518);
  not NOT_2743(g9976,g2537);
  not NOT_2744(g9977,g2667);
  not NOT_2745(g9978,g2756);
  not NOT_2746(g9982,g3976);
  not NOT_2747(g9983,g4239);
  not NOT_2748(g9985,g4332);
  not NOT_2749(g9989,g5077);
  not NOT_2750(g9992,g5990);
  not NOT_2751(g9995,g6035);
  not NOT_2752(g9999,g6109);
  not NOT_2753(g10000,g6151);
  not NOT_2754(g10001,g6105);
  not NOT_2755(g10002,g6195);
  not NOT_2756(I13539,g6381);
  not NOT_2757(g10003,I13539);
  not NOT_2758(g10014,g6439);
  not NOT_2759(g10019,g6479);
  not NOT_2760(g10026,g6494);
  not NOT_2761(g10027,g6523);
  not NOT_2762(g10028,g8);
  not NOT_2763(I13548,g94);
  not NOT_2764(g10029,I13548);
  not NOT_2765(g10030,g116);
  not NOT_2766(I13552,g121);
  not NOT_2767(g10031,I13552);
  not NOT_2768(g10032,g562);
  not NOT_2769(g10033,g655);
  not NOT_2770(g10035,g1720);
  not NOT_2771(g10036,g1816);
  not NOT_2772(g10037,g1848);
  not NOT_2773(g10038,g2241);
  not NOT_2774(g10039,g2273);
  not NOT_2775(g10040,g2652);
  not NOT_2776(g10042,g2671);
  not NOT_2777(g10043,g1632);
  not NOT_2778(g10044,g5357);
  not NOT_2779(g10047,g5421);
  not NOT_2780(g10050,g6336);
  not NOT_2781(g10053,g6381);
  not NOT_2782(g10057,g6455);
  not NOT_2783(g10058,g6497);
  not NOT_2784(g10059,g6451);
  not NOT_2785(g10060,g6541);
  not NOT_2786(I13581,g6727);
  not NOT_2787(g10061,I13581);
  not NOT_2788(g10072,g9);
  not NOT_2789(g10073,g134);
  not NOT_2790(g10074,g718);
  not NOT_2791(g10077,g1724);
  not NOT_2792(g10078,g1854);
  not NOT_2793(g10079,g1950);
  not NOT_2794(g10080,g1982);
  not NOT_2795(g10081,g2279);
  not NOT_2796(g10082,g2375);
  not NOT_2797(g10083,g2407);
  not NOT_2798(g10084,g2837);
  not NOT_2799(g10085,g1768);
  not NOT_2800(g10086,g2193);
  not NOT_2801(I13597,g4417);
  not NOT_2802(g10087,I13597);
  not NOT_2803(g10090,g5348);
  not NOT_2804(g10093,g5703);
  not NOT_2805(g10096,g5767);
  not NOT_2806(g10099,g6682);
  not NOT_2807(g10102,g6727);
  not NOT_2808(g10106,g16);
  not NOT_2809(I13606,g74);
  not NOT_2810(g10107,I13606);
  not NOT_2811(g10108,g120);
  not NOT_2812(g10109,g135);
  not NOT_2813(g10110,g661);
  not NOT_2814(g10111,g1858);
  not NOT_2815(g10112,g1988);
  not NOT_2816(g10113,g2084);
  not NOT_2817(g10114,g2116);
  not NOT_2818(g10115,g2283);
  not NOT_2819(g10116,g2413);
  not NOT_2820(g10117,g2509);
  not NOT_2821(g10118,g2541);
  not NOT_2822(g10119,g2841);
  not NOT_2823(g10120,g1902);
  not NOT_2824(g10121,g2327);
  not NOT_2825(I13623,g4294);
  not NOT_2826(g10122,I13623);
  not NOT_2827(g10129,g5352);
  not NOT_2828(g10130,g5694);
  not NOT_2829(g10133,g6049);
  not NOT_2830(g10136,g6113);
  not NOT_2831(g10139,g136);
  not NOT_2832(g10140,g19);
  not NOT_2833(I13634,g79);
  not NOT_2834(g10141,I13634);
  not NOT_2835(I13637,g102);
  not NOT_2836(g10142,I13637);
  not NOT_2837(g10143,g568);
  not NOT_2838(g10147,g728);
  not NOT_2839(g10150,g1700);
  not NOT_2840(g10151,g1992);
  not NOT_2841(g10152,g2122);
  not NOT_2842(g10153,g2417);
  not NOT_2843(g10154,g2547);
  not NOT_2844(g10155,g2643);
  not NOT_2845(g10156,g2675);
  not NOT_2846(g10157,g2036);
  not NOT_2847(g10158,g2461);
  not NOT_2848(g10159,g4477);
  not NOT_2849(g10165,g5698);
  not NOT_2850(g10166,g6040);
  not NOT_2851(g10169,g6395);
  not NOT_2852(g10172,g6459);
  not NOT_2853(g10175,g28);
  not NOT_2854(g10176,g44);
  not NOT_2855(g10177,g1834);
  not NOT_2856(g10178,g2126);
  not NOT_2857(g10180,g2259);
  not NOT_2858(g10181,g2551);
  not NOT_2859(g10182,g2681);
  not NOT_2860(g10183,g2595);
  not NOT_2861(g10184,g4486);
  not NOT_2862(g10190,g6044);
  not NOT_2863(g10191,g6386);
  not NOT_2864(g10194,g6741);
  not NOT_2865(g10197,g31);
  not NOT_2866(I13672,g106);
  not NOT_2867(g10198,I13672);
  not NOT_2868(g10199,g1968);
  not NOT_2869(g10200,g2138);
  not NOT_2870(g10203,g2393);
  not NOT_2871(g10204,g2685);
  not NOT_2872(g10206,g4489);
  not NOT_2873(g10212,g6390);
  not NOT_2874(g10213,g6732);
  not NOT_2875(I13684,g128);
  not NOT_2876(g10216,I13684);
  not NOT_2877(g10217,g2102);
  not NOT_2878(g10218,g2527);
  not NOT_2879(g10219,g2697);
  not NOT_2880(g10222,g4492);
  not NOT_2881(g10223,g4561);
  not NOT_2882(g10229,g6736);
  not NOT_2883(I13694,g117);
  not NOT_2884(g10230,I13694);
  not NOT_2885(g10231,g2661);
  not NOT_2886(g10232,g4527);
  not NOT_2887(I13699,g4581);
  not NOT_2888(g10233,I13699);
  not NOT_2889(g10261,g4555);
  not NOT_2890(g10262,g586);
  not NOT_2891(I13705,g63);
  not NOT_2892(g10272,I13705);
  not NOT_2893(I13708,g136);
  not NOT_2894(g10273,I13708);
  not NOT_2895(g10274,g976);
  not NOT_2896(g10275,g4584);
  not NOT_2897(g10278,g4628);
  not NOT_2898(I13715,g71);
  not NOT_2899(g10287,I13715);
  not NOT_2900(I13718,g890);
  not NOT_2901(g10288,I13718);
  not NOT_2902(g10289,g1319);
  not NOT_2903(I13723,g3167);
  not NOT_2904(g10295,I13723);
  not NOT_2905(I13726,g4537);
  not NOT_2906(g10306,I13726);
  not NOT_2907(g10308,g4459);
  not NOT_2908(g10311,g4633);
  not NOT_2909(I13740,g85);
  not NOT_2910(g10319,I13740);
  not NOT_2911(g10320,g817);
  not NOT_2912(I13744,g3518);
  not NOT_2913(g10323,I13744);
  not NOT_2914(g10334,g4420);
  not NOT_2915(g10335,g4483);
  not NOT_2916(g10337,g5016);
  not NOT_2917(I13759,g6754);
  not NOT_2918(g10347,I13759);
  not NOT_2919(I13762,g6755);
  not NOT_2920(g10348,I13762);
  not NOT_2921(g10349,g6956);
  not NOT_2922(g10350,g6800);
  not NOT_2923(g10351,g6802);
  not NOT_2924(g10352,g6804);
  not NOT_2925(g10353,g6803);
  not NOT_2926(g10354,g6811);
  not NOT_2927(g10355,g6816);
  not NOT_2928(g10356,g6819);
  not NOT_2929(g10357,g6825);
  not NOT_2930(g10358,g6827);
  not NOT_2931(g10359,g6830);
  not NOT_2932(g10360,g6836);
  not NOT_2933(g10361,g6841);
  not NOT_2934(g10362,g6850);
  not NOT_2935(I13779,g6868);
  not NOT_2936(g10363,I13779);
  not NOT_2937(g10364,g6869);
  not NOT_2938(g10365,g6867);
  not NOT_2939(g10366,g6895);
  not NOT_2940(g10367,g6870);
  not NOT_2941(g10368,g6887);
  not NOT_2942(g10369,g6873);
  not NOT_2943(g10370,g7095);
  not NOT_2944(g10371,g6918);
  not NOT_2945(g10372,g6900);
  not NOT_2946(g10373,g6917);
  not NOT_2947(g10374,g6903);
  not NOT_2948(g10375,g6941);
  not NOT_2949(g10376,g6923);
  not NOT_2950(g10377,g6940);
  not NOT_2951(g10378,g6926);
  not NOT_2952(g10379,g6953);
  not NOT_2953(g10380,g6960);
  not NOT_2954(g10381,g6957);
  not NOT_2955(g10382,g6958);
  not NOT_2956(g10383,g6978);
  not NOT_2957(I13802,g6971);
  not NOT_2958(g10384,I13802);
  not NOT_2959(I13805,g6976);
  not NOT_2960(g10385,I13805);
  not NOT_2961(g10386,g6982);
  not NOT_2962(g10387,g6996);
  not NOT_2963(g10388,g6983);
  not NOT_2964(g10389,g6986);
  not NOT_2965(g10390,g6987);
  not NOT_2966(g10391,g6988);
  not NOT_2967(g10392,g6989);
  not NOT_2968(g10393,g6991);
  not NOT_2969(g10394,g6994);
  not NOT_2970(g10395,g6995);
  not NOT_2971(g10396,g6997);
  not NOT_2972(g10397,g7018);
  not NOT_2973(g10398,g6999);
  not NOT_2974(g10399,g7017);
  not NOT_2975(g10400,g7002);
  not NOT_2976(g10401,g7041);
  not NOT_2977(g10402,g7023);
  not NOT_2978(g10403,g7040);
  not NOT_2979(g10404,g7026);
  not NOT_2980(g10405,g7064);
  not NOT_2981(g10406,g7046);
  not NOT_2982(g10407,g7063);
  not NOT_2983(g10408,g7049);
  not NOT_2984(g10409,g7087);
  not NOT_2985(g10410,g7069);
  not NOT_2986(g10411,g7086);
  not NOT_2987(g10412,g7072);
  not NOT_2988(g10413,g7110);
  not NOT_2989(g10414,g7092);
  not NOT_2990(g10415,g7109);
  not NOT_2991(g10416,g10318);
  not NOT_2992(g10417,g7117);
  not NOT_2993(g10418,g8818);
  not NOT_2994(g10419,g8821);
  not NOT_2995(g10420,g9239);
  not NOT_2996(g10427,g10053);
  not NOT_2997(g10428,g9631);
  not NOT_2998(g10429,g7148);
  not NOT_2999(I13847,g7266);
  not NOT_3000(g10430,I13847);
  not NOT_3001(I13857,g9780);
  not NOT_3002(g10473,I13857);
  not NOT_3003(g10474,g8841);
  not NOT_3004(g10475,g8844);
  not NOT_3005(g10487,g10233);
  not NOT_3006(g10489,g9259);
  not NOT_3007(g10490,g9274);
  not NOT_3008(g10497,g10102);
  not NOT_3009(g10498,g7161);
  not NOT_3010(I13872,g7474);
  not NOT_3011(g10499,I13872);
  not NOT_3012(I13875,g1233);
  not NOT_3013(g10500,I13875);
  not NOT_3014(g10502,g8876);
  not NOT_3015(g10503,g8879);
  not NOT_3016(g10504,g8763);
  not NOT_3017(g10509,g10233);
  not NOT_3018(g10518,g9311);
  not NOT_3019(g10519,g9326);
  not NOT_3020(I13889,g7598);
  not NOT_3021(g10521,I13889);
  not NOT_3022(I13892,g1576);
  not NOT_3023(g10527,I13892);
  not NOT_3024(g10530,g8922);
  not NOT_3025(g10531,g8925);
  not NOT_3026(g10532,g10233);
  not NOT_3027(g10533,g8795);
  not NOT_3028(g10540,g9392);
  not NOT_3029(g10541,g9407);
  not NOT_3030(g10542,g7196);
  not NOT_3031(I13906,g7620);
  not NOT_3032(g10544,I13906);
  not NOT_3033(g10553,g8971);
  not NOT_3034(g10554,g8974);
  not NOT_3035(g10564,g9462);
  not NOT_3036(g10570,g9021);
  not NOT_3037(g10571,g10233);
  not NOT_3038(g10572,g10233);
  not NOT_3039(g10581,g9529);
  not NOT_3040(g10582,g7116);
  not NOT_3041(g10597,g10233);
  not NOT_3042(g10606,g10233);
  not NOT_3043(g10607,g10233);
  not NOT_3044(g10608,g9155);
  not NOT_3045(g10612,g10233);
  not NOT_3046(g10613,g10233);
  not NOT_3047(g10620,g10233);
  not NOT_3048(g10621,g7567);
  not NOT_3049(I13968,g7697);
  not NOT_3050(g10627,I13968);
  not NOT_3051(g10652,g7601);
  not NOT_3052(I13979,g7733);
  not NOT_3053(g10658,I13979);
  not NOT_3054(g10664,g8928);
  not NOT_3055(I13990,g7636);
  not NOT_3056(g10678,I13990);
  not NOT_3057(I13995,g8744);
  not NOT_3058(g10685,I13995);
  not NOT_3059(g10708,g7836);
  not NOT_3060(I14006,g9104);
  not NOT_3061(g10710,I14006);
  not NOT_3062(g10725,g7846);
  not NOT_3063(I14016,g9104);
  not NOT_3064(g10727,I14016);
  not NOT_3065(g10741,g8411);
  not NOT_3066(g10761,g8411);
  not NOT_3067(g10762,g8470);
  not NOT_3068(I14033,g8912);
  not NOT_3069(g10776,I14033);
  not NOT_3070(g10794,g8470);
  not NOT_3071(g10795,g7202);
  not NOT_3072(g10804,g9772);
  not NOT_3073(I14046,g9900);
  not NOT_3074(g10805,I14046);
  not NOT_3075(I14050,g9963);
  not NOT_3076(g10812,I14050);
  not NOT_3077(g10815,g9917);
  not NOT_3078(I14054,g10028);
  not NOT_3079(g10816,I14054);
  not NOT_3080(g10830,g10087);
  not NOT_3081(I14069,g9104);
  not NOT_3082(g10851,I14069);
  not NOT_3083(g10857,g8712);
  not NOT_3084(g10872,g7567);
  not NOT_3085(I14079,g7231);
  not NOT_3086(g10877,I14079);
  not NOT_3087(g10881,g7567);
  not NOT_3088(g10882,g7601);
  not NOT_3089(g10897,g7601);
  not NOT_3090(g10960,g9007);
  not NOT_3091(g10980,g9051);
  not NOT_3092(I14119,g7824);
  not NOT_3093(g10981,I14119);
  not NOT_3094(g11011,g10274);
  not NOT_3095(g11017,g10289);
  not NOT_3096(g11026,g8434);
  not NOT_3097(g11030,g8292);
  not NOT_3098(g11031,g8609);
  not NOT_3099(g11033,g8500);
  not NOT_3100(g11034,g7611);
  not NOT_3101(g11038,g8632);
  not NOT_3102(g11042,g8691);
  not NOT_3103(g11043,g8561);
  not NOT_3104(I14158,g8806);
  not NOT_3105(g11048,I14158);
  not NOT_3106(g11110,g8728);
  not NOT_3107(g11122,g8751);
  not NOT_3108(g11128,g7993);
  not NOT_3109(g11129,g7994);
  not NOT_3110(I14192,g10233);
  not NOT_3111(g11136,I14192);
  not NOT_3112(g11143,g8032);
  not NOT_3113(g11147,g8417);
  not NOT_3114(g11164,g8085);
  not NOT_3115(I14222,g8286);
  not NOT_3116(g11165,I14222);
  not NOT_3117(g11170,g8476);
  not NOT_3118(g11181,g8134);
  not NOT_3119(I14241,g8356);
  not NOT_3120(g11182,I14241);
  not NOT_3121(g11183,g8135);
  not NOT_3122(g11192,g8038);
  not NOT_3123(I14267,g7835);
  not NOT_3124(g11202,I14267);
  not NOT_3125(I14271,g8456);
  not NOT_3126(g11204,I14271);
  not NOT_3127(g11214,g9602);
  not NOT_3128(g11215,g8285);
  not NOT_3129(g11233,g9664);
  not NOT_3130(g11234,g8355);
  not NOT_3131(I14301,g8571);
  not NOT_3132(g11235,I14301);
  not NOT_3133(g11236,g8357);
  not NOT_3134(I14305,g8805);
  not NOT_3135(g11237,I14305);
  not NOT_3136(g11249,g8405);
  not NOT_3137(g11250,g7502);
  not NOT_3138(g11268,g7515);
  not NOT_3139(g11269,g7516);
  not NOT_3140(I14326,g8607);
  not NOT_3141(g11290,I14326);
  not NOT_3142(g11291,g7526);
  not NOT_3143(g11293,g7527);
  not NOT_3144(g11294,g7598);
  not NOT_3145(g11316,g8967);
  not NOT_3146(I14346,g10233);
  not NOT_3147(g11317,I14346);
  not NOT_3148(g11324,g7542);
  not NOT_3149(g11325,g7543);
  not NOT_3150(g11336,g7620);
  not NOT_3151(g11344,g9015);
  not NOT_3152(I14365,g3303);
  not NOT_3153(g11349,I14365);
  not NOT_3154(I14381,g8300);
  not NOT_3155(g11367,I14381);
  not NOT_3156(g11371,g7565);
  not NOT_3157(g11373,g7566);
  not NOT_3158(g11383,g9061);
  not NOT_3159(I14395,g3654);
  not NOT_3160(g11388,I14395);
  not NOT_3161(I14409,g8364);
  not NOT_3162(g11398,I14409);
  not NOT_3163(g11401,g7593);
  not NOT_3164(g11402,g7594);
  not NOT_3165(g11403,g7595);
  not NOT_3166(g11404,g7596);
  not NOT_3167(g11413,g9100);
  not NOT_3168(I14424,g4005);
  not NOT_3169(g11418,I14424);
  not NOT_3170(g11425,g7640);
  not NOT_3171(g11428,g7615);
  not NOT_3172(g11429,g7616);
  not NOT_3173(g11430,g7617);
  not NOT_3174(g11431,g7618);
  not NOT_3175(I14450,g4191);
  not NOT_3176(g11447,I14450);
  not NOT_3177(I14455,g10197);
  not NOT_3178(g11450,I14455);
  not NOT_3179(g11467,g7623);
  not NOT_3180(g11468,g7624);
  not NOT_3181(g11470,g7625);
  not NOT_3182(g11471,g7626);
  not NOT_3183(g11472,g7918);
  not NOT_3184(I14475,g10175);
  not NOT_3185(g11498,I14475);
  not NOT_3186(g11509,g7632);
  not NOT_3187(g11510,g7633);
  not NOT_3188(g11512,g7634);
  not NOT_3189(g11513,g7948);
  not NOT_3190(g11519,g8481);
  not NOT_3191(I14505,g10140);
  not NOT_3192(g11547,I14505);
  not NOT_3193(g11560,g7647);
  not NOT_3194(g11562,g7648);
  not NOT_3195(g11576,g8542);
  not NOT_3196(I14537,g10106);
  not NOT_3197(g11592,I14537);
  not NOT_3198(g11608,g7659);
  not NOT_3199(g11609,g7660);
  not NOT_3200(g11615,g6875);
  not NOT_3201(g11631,g8595);
  not NOT_3202(I14550,g10072);
  not NOT_3203(g11640,I14550);
  not NOT_3204(g11652,g7674);
  not NOT_3205(g11663,g6905);
  not NOT_3206(g11677,g7689);
  not NOT_3207(I14563,g802);
  not NOT_3208(g11678,I14563);
  not NOT_3209(I14567,g9708);
  not NOT_3210(g11686,I14567);
  not NOT_3211(I14570,g7932);
  not NOT_3212(g11691,I14570);
  not NOT_3213(g11702,g6928);
  not NOT_3214(I14576,g8791);
  not NOT_3215(g11705,I14576);
  not NOT_3216(I14579,g8792);
  not NOT_3217(g11706,I14579);
  not NOT_3218(I14584,g9766);
  not NOT_3219(g11709,I14584);
  not NOT_3220(g11714,g8107);
  not NOT_3221(I14589,g8818);
  not NOT_3222(g11720,I14589);
  not NOT_3223(g11721,g10074);
  not NOT_3224(I14593,g9978);
  not NOT_3225(g11724,I14593);
  not NOT_3226(g11735,g8534);
  not NOT_3227(g11736,g8165);
  not NOT_3228(g11741,g10033);
  not NOT_3229(I14602,g9340);
  not NOT_3230(g11744,I14602);
  not NOT_3231(g11753,g8587);
  not NOT_3232(g11754,g8229);
  not NOT_3233(g11762,g7964);
  not NOT_3234(g11769,g8626);
  not NOT_3235(I14619,g4185);
  not NOT_3236(g11770,I14619);
  not NOT_3237(I14623,g8925);
  not NOT_3238(g11772,I14623);
  not NOT_3239(g11779,g9602);
  not NOT_3240(g11786,g7549);
  not NOT_3241(I14630,g7717);
  not NOT_3242(g11790,I14630);
  not NOT_3243(I14633,g9340);
  not NOT_3244(g11793,I14633);
  not NOT_3245(g11796,g7985);
  not NOT_3246(g11810,g9664);
  not NOT_3247(g11811,g9724);
  not NOT_3248(g11812,g7567);
  not NOT_3249(g11815,g7582);
  not NOT_3250(g11819,g7717);
  not NOT_3251(I14644,g7717);
  not NOT_3252(g11820,I14644);
  not NOT_3253(I14647,g7717);
  not NOT_3254(g11823,I14647);
  not NOT_3255(I14650,g9340);
  not NOT_3256(g11826,I14650);
  not NOT_3257(I14653,g9417);
  not NOT_3258(g11829,I14653);
  not NOT_3259(g11832,g8011);
  not NOT_3260(g11833,g8026);
  not NOT_3261(g11841,g9800);
  not NOT_3262(I14660,g9746);
  not NOT_3263(g11842,I14660);
  not NOT_3264(I14663,g9747);
  not NOT_3265(g11845,I14663);
  not NOT_3266(g11849,g7601);
  not NOT_3267(I14668,g7753);
  not NOT_3268(g11852,I14668);
  not NOT_3269(I14671,g7717);
  not NOT_3270(g11855,I14671);
  not NOT_3271(g11861,g8070);
  not NOT_3272(g11865,g10124);
  not NOT_3273(g11866,g9883);
  not NOT_3274(I14679,g9332);
  not NOT_3275(g11867,I14679);
  not NOT_3276(g11868,g9185);
  not NOT_3277(I14684,g7717);
  not NOT_3278(g11872,I14684);
  not NOT_3279(I14687,g7753);
  not NOT_3280(g11875,I14687);
  not NOT_3281(I14690,g9340);
  not NOT_3282(g11878,I14690);
  not NOT_3283(g11884,g8125);
  not NOT_3284(g11888,g10160);
  not NOT_3285(g11889,g9954);
  not NOT_3286(I14702,g7717);
  not NOT_3287(g11894,I14702);
  not NOT_3288(I14705,g7717);
  not NOT_3289(g11897,I14705);
  not NOT_3290(I14708,g9417);
  not NOT_3291(g11900,I14708);
  not NOT_3292(g11910,g10185);
  not NOT_3293(g11911,g10022);
  not NOT_3294(g11912,g8989);
  not NOT_3295(I14727,g7753);
  not NOT_3296(g11917,I14727);
  not NOT_3297(I14730,g7717);
  not NOT_3298(g11920,I14730);
  not NOT_3299(g11927,g10207);
  not NOT_3300(I14742,g9534);
  not NOT_3301(g11928,I14742);
  not NOT_3302(I14745,g10029);
  not NOT_3303(g11929,I14745);
  not NOT_3304(g11930,g9281);
  not NOT_3305(I14749,g10031);
  not NOT_3306(g11931,I14749);
  not NOT_3307(I14761,g7753);
  not NOT_3308(g11941,I14761);
  not NOT_3309(g11948,g10224);
  not NOT_3310(I14773,g9581);
  not NOT_3311(g11949,I14773);
  not NOT_3312(g11963,g9153);
  not NOT_3313(g11964,g9154);
  not NOT_3314(I14797,g9636);
  not NOT_3315(g11965,I14797);
  not NOT_3316(I14800,g10107);
  not NOT_3317(g11966,I14800);
  not NOT_3318(I14823,g8056);
  not NOT_3319(g11981,I14823);
  not NOT_3320(g11984,g9186);
  not NOT_3321(I14827,g9686);
  not NOT_3322(g11985,I14827);
  not NOT_3323(I14830,g10141);
  not NOT_3324(g11986,I14830);
  not NOT_3325(I14833,g10142);
  not NOT_3326(g11987,I14833);
  not NOT_3327(I14836,g9688);
  not NOT_3328(g11988,I14836);
  not NOT_3329(I14839,g9689);
  not NOT_3330(g11989,I14839);
  not NOT_3331(g11991,g9485);
  not NOT_3332(I14862,g8092);
  not NOT_3333(g12009,I14862);
  not NOT_3334(g12012,g9213);
  not NOT_3335(I14866,g9748);
  not NOT_3336(g12013,I14866);
  not NOT_3337(g12018,g9538);
  not NOT_3338(g12021,g9543);
  not NOT_3339(g12036,g9245);
  not NOT_3340(I14893,g9819);
  not NOT_3341(g12037,I14893);
  not NOT_3342(I14896,g9820);
  not NOT_3343(g12038,I14896);
  not NOT_3344(I14899,g10198);
  not NOT_3345(g12039,I14899);
  not NOT_3346(I14902,g9821);
  not NOT_3347(g12040,I14902);
  not NOT_3348(I14905,g9822);
  not NOT_3349(g12041,I14905);
  not NOT_3350(g12047,g9591);
  not NOT_3351(g12051,g9595);
  not NOT_3352(g12054,g7690);
  not NOT_3353(I14932,g9901);
  not NOT_3354(g12074,I14932);
  not NOT_3355(I14935,g9902);
  not NOT_3356(g12075,I14935);
  not NOT_3357(g12076,g9280);
  not NOT_3358(I14939,g10216);
  not NOT_3359(g12077,I14939);
  not NOT_3360(g12082,g9645);
  not NOT_3361(g12086,g9654);
  not NOT_3362(g12088,g7701);
  not NOT_3363(g12107,g9687);
  not NOT_3364(I14964,g10230);
  not NOT_3365(g12108,I14964);
  not NOT_3366(I14967,g9964);
  not NOT_3367(g12109,I14967);
  not NOT_3368(I14970,g9965);
  not NOT_3369(g12110,I14970);
  not NOT_3370(g12122,g9705);
  not NOT_3371(I14999,g10030);
  not NOT_3372(g12143,I14999);
  not NOT_3373(g12180,g9477);
  not NOT_3374(g12181,g9478);
  not NOT_3375(I15030,g10073);
  not NOT_3376(g12182,I15030);
  not NOT_3377(I15033,g10273);
  not NOT_3378(g12183,I15033);
  not NOT_3379(I15036,g799);
  not NOT_3380(g12184,I15036);
  not NOT_3381(I15070,g10108);
  not NOT_3382(g12217,I15070);
  not NOT_3383(I15073,g10109);
  not NOT_3384(g12218,I15073);
  not NOT_3385(g12233,g10338);
  not NOT_3386(I15102,g5313);
  not NOT_3387(g12238,I15102);
  not NOT_3388(g12295,g7139);
  not NOT_3389(I15144,g5659);
  not NOT_3390(g12300,I15144);
  not NOT_3391(g12321,g9637);
  not NOT_3392(I15162,g10176);
  not NOT_3393(g12322,I15162);
  not NOT_3394(g12337,g9340);
  not NOT_3395(g12345,g7158);
  not NOT_3396(I15190,g6005);
  not NOT_3397(g12350,I15190);
  not NOT_3398(I15205,g10139);
  not NOT_3399(g12367,I15205);
  not NOT_3400(I15208,g637);
  not NOT_3401(g12368,I15208);
  not NOT_3402(g12378,g9417);
  not NOT_3403(I15223,g10119);
  not NOT_3404(g12381,I15223);
  not NOT_3405(g12399,g9920);
  not NOT_3406(g12417,g7175);
  not NOT_3407(I15238,g6351);
  not NOT_3408(g12422,I15238);
  not NOT_3409(I15250,g9152);
  not NOT_3410(g12430,I15250);
  not NOT_3411(g12440,g9985);
  not NOT_3412(g12465,g7192);
  not NOT_3413(I15284,g6697);
  not NOT_3414(g12470,I15284);
  not NOT_3415(I15295,g8515);
  not NOT_3416(g12477,I15295);
  not NOT_3417(g12487,g9340);
  not NOT_3418(I15316,g10087);
  not NOT_3419(g12490,I15316);
  not NOT_3420(g12497,g9780);
  not NOT_3421(g12543,g9417);
  not NOT_3422(g12546,g8740);
  not NOT_3423(g12563,g9864);
  not NOT_3424(g12598,g7004);
  not NOT_3425(g12614,g9935);
  not NOT_3426(I15382,g9071);
  not NOT_3427(g12640,I15382);
  not NOT_3428(g12656,g7028);
  not NOT_3429(g12672,g10003);
  not NOT_3430(g12705,g7051);
  not NOT_3431(g12721,g10061);
  not NOT_3432(g12738,g9374);
  not NOT_3433(g12749,g7074);
  not NOT_3434(g12760,g10272);
  not NOT_3435(g12778,g9856);
  not NOT_3436(g12779,g9444);
  not NOT_3437(g12790,g7097);
  not NOT_3438(g12793,g10287);
  not NOT_3439(g12804,g9927);
  not NOT_3440(g12805,g9511);
  not NOT_3441(g12811,g10319);
  not NOT_3442(g12818,g8792);
  not NOT_3443(g12820,g10233);
  not NOT_3444(g12823,g9206);
  not NOT_3445(g12830,g9995);
  not NOT_3446(g12831,g9569);
  not NOT_3447(I15448,g10877);
  not NOT_3448(g12833,I15448);
  not NOT_3449(g12834,g10349);
  not NOT_3450(g12835,g10352);
  not NOT_3451(g12836,g10351);
  not NOT_3452(g12837,g10354);
  not NOT_3453(g12838,g10353);
  not NOT_3454(g12839,g10350);
  not NOT_3455(g12840,g10356);
  not NOT_3456(g12841,g10357);
  not NOT_3457(g12842,g10355);
  not NOT_3458(g12843,g10359);
  not NOT_3459(g12844,g10360);
  not NOT_3460(g12845,g10358);
  not NOT_3461(I15474,g10364);
  not NOT_3462(g12857,I15474);
  not NOT_3463(g12859,g10366);
  not NOT_3464(g12860,g10368);
  not NOT_3465(g12861,g10367);
  not NOT_3466(g12862,g10370);
  not NOT_3467(g12863,g10371);
  not NOT_3468(g12864,g10373);
  not NOT_3469(g12865,g10372);
  not NOT_3470(g12866,g10369);
  not NOT_3471(g12867,g10375);
  not NOT_3472(g12868,g10377);
  not NOT_3473(g12869,g10376);
  not NOT_3474(g12870,g10374);
  not NOT_3475(g12871,g10378);
  not NOT_3476(g12872,g10379);
  not NOT_3477(g12873,g10380);
  not NOT_3478(g12874,g10383);
  not NOT_3479(I15494,g10385);
  not NOT_3480(g12875,I15494);
  not NOT_3481(g12878,g10386);
  not NOT_3482(g12879,g10381);
  not NOT_3483(g12880,g10387);
  not NOT_3484(g12881,g10388);
  not NOT_3485(g12882,g10389);
  not NOT_3486(g12883,g10390);
  not NOT_3487(g12884,g10392);
  not NOT_3488(g12885,g10382);
  not NOT_3489(g12886,g10393);
  not NOT_3490(g12887,g10394);
  not NOT_3491(g12888,g10395);
  not NOT_3492(g12889,g10396);
  not NOT_3493(g12890,g10397);
  not NOT_3494(g12891,g10399);
  not NOT_3495(g12892,g10398);
  not NOT_3496(g12893,g10391);
  not NOT_3497(g12894,g10401);
  not NOT_3498(g12895,g10403);
  not NOT_3499(g12896,g10402);
  not NOT_3500(g12897,g10400);
  not NOT_3501(g12898,g10405);
  not NOT_3502(g12899,g10407);
  not NOT_3503(g12900,g10406);
  not NOT_3504(g12901,g10404);
  not NOT_3505(g12902,g10409);
  not NOT_3506(g12903,g10411);
  not NOT_3507(g12904,g10410);
  not NOT_3508(g12905,g10408);
  not NOT_3509(g12906,g10413);
  not NOT_3510(g12907,g10415);
  not NOT_3511(g12908,g10414);
  not NOT_3512(g12909,g10412);
  not NOT_3513(g12914,g12235);
  not NOT_3514(I15533,g11867);
  not NOT_3515(g12918,I15533);
  not NOT_3516(I15536,g1227);
  not NOT_3517(g12919,I15536);
  not NOT_3518(g12921,g12228);
  not NOT_3519(g12922,g12297);
  not NOT_3520(I15542,g1570);
  not NOT_3521(g12923,I15542);
  not NOT_3522(g12929,g12550);
  not NOT_3523(g12930,g12347);
  not NOT_3524(I15550,g10430);
  not NOT_3525(g12932,I15550);
  not NOT_3526(g12936,g12601);
  not NOT_3527(g12937,g12419);
  not NOT_3528(I15556,g11928);
  not NOT_3529(g12938,I15556);
  not NOT_3530(g12940,g11744);
  not NOT_3531(g12944,g12659);
  not NOT_3532(g12945,g12467);
  not NOT_3533(I15564,g11949);
  not NOT_3534(g12946,I15564);
  not NOT_3535(g12950,g12708);
  not NOT_3536(I15569,g11965);
  not NOT_3537(g12951,I15569);
  not NOT_3538(I15572,g10499);
  not NOT_3539(g12952,I15572);
  not NOT_3540(I15577,g10430);
  not NOT_3541(g12955,I15577);
  not NOT_3542(g12967,g11790);
  not NOT_3543(g12968,g11793);
  not NOT_3544(g12975,g12752);
  not NOT_3545(I15587,g11985);
  not NOT_3546(g12976,I15587);
  not NOT_3547(I15590,g11988);
  not NOT_3548(g12977,I15590);
  not NOT_3549(I15593,g11989);
  not NOT_3550(g12978,I15593);
  not NOT_3551(I15600,g10430);
  not NOT_3552(g12983,I15600);
  not NOT_3553(g12995,g11820);
  not NOT_3554(g12996,g11823);
  not NOT_3555(g12997,g11826);
  not NOT_3556(g12998,g11829);
  not NOT_3557(I15609,g12013);
  not NOT_3558(g13003,I15609);
  not NOT_3559(g13007,g11852);
  not NOT_3560(g13008,g11855);
  not NOT_3561(I15617,g12037);
  not NOT_3562(g13009,I15617);
  not NOT_3563(I15620,g12038);
  not NOT_3564(g13010,I15620);
  not NOT_3565(I15623,g12040);
  not NOT_3566(g13011,I15623);
  not NOT_3567(I15626,g12041);
  not NOT_3568(g13012,I15626);
  not NOT_3569(g13014,g11872);
  not NOT_3570(g13015,g11875);
  not NOT_3571(g13016,g11878);
  not NOT_3572(I15633,g12074);
  not NOT_3573(g13017,I15633);
  not NOT_3574(I15636,g12075);
  not NOT_3575(g13018,I15636);
  not NOT_3576(g13022,g11894);
  not NOT_3577(g13023,g11897);
  not NOT_3578(g13024,g11900);
  not NOT_3579(g13026,g11018);
  not NOT_3580(I15647,g12109);
  not NOT_3581(g13027,I15647);
  not NOT_3582(I15650,g12110);
  not NOT_3583(g13028,I15650);
  not NOT_3584(g13033,g11917);
  not NOT_3585(g13034,g11920);
  not NOT_3586(g13036,g10981);
  not NOT_3587(g13037,g10981);
  not NOT_3588(I15663,g5308);
  not NOT_3589(g13039,I15663);
  not NOT_3590(I15667,g12143);
  not NOT_3591(g13041,I15667);
  not NOT_3592(g13045,g11941);
  not NOT_3593(I15677,g5654);
  not NOT_3594(g13049,I15677);
  not NOT_3595(g13051,g11964);
  not NOT_3596(I15682,g12182);
  not NOT_3597(g13055,I15682);
  not NOT_3598(g13061,g10981);
  not NOT_3599(g13062,g10981);
  not NOT_3600(g13064,g11705);
  not NOT_3601(g13065,g10476);
  not NOT_3602(I15697,g6000);
  not NOT_3603(g13068,I15697);
  not NOT_3604(g13070,g11984);
  not NOT_3605(I15702,g12217);
  not NOT_3606(g13074,I15702);
  not NOT_3607(I15705,g12218);
  not NOT_3608(g13075,I15705);
  not NOT_3609(g13082,g10981);
  not NOT_3610(I15717,g6346);
  not NOT_3611(g13085,I15717);
  not NOT_3612(g13087,g12012);
  not NOT_3613(I15727,g10981);
  not NOT_3614(g13096,I15727);
  not NOT_3615(I15732,g6692);
  not NOT_3616(g13099,I15732);
  not NOT_3617(I15736,g12322);
  not NOT_3618(g13101,I15736);
  not NOT_3619(g13103,g10905);
  not NOT_3620(g13106,g10981);
  not NOT_3621(g13107,g10476);
  not NOT_3622(g13116,g10935);
  not NOT_3623(g13117,g10981);
  not NOT_3624(g13120,g10632);
  not NOT_3625(g13132,g10632);
  not NOT_3626(g13133,g11330);
  not NOT_3627(I15765,g10823);
  not NOT_3628(g13138,I15765);
  not NOT_3629(g13140,g10632);
  not NOT_3630(g13141,g11374);
  not NOT_3631(g13142,g10632);
  not NOT_3632(I15773,g10430);
  not NOT_3633(g13144,I15773);
  not NOT_3634(g13173,g10632);
  not NOT_3635(g13174,g10741);
  not NOT_3636(g13175,g10909);
  not NOT_3637(I15782,g10430);
  not NOT_3638(g13177,I15782);
  not NOT_3639(g13188,g10909);
  not NOT_3640(g13189,g10762);
  not NOT_3641(g13190,g10939);
  not NOT_3642(I15788,g10430);
  not NOT_3643(g13191,I15788);
  not NOT_3644(g13209,g10632);
  not NOT_3645(g13215,g10909);
  not NOT_3646(g13216,g10939);
  not NOT_3647(g13222,g10590);
  not NOT_3648(I15800,g11607);
  not NOT_3649(g13223,I15800);
  not NOT_3650(g13239,g10632);
  not NOT_3651(g13246,g10939);
  not NOT_3652(g13249,g10590);
  not NOT_3653(I15811,g11128);
  not NOT_3654(g13250,I15811);
  not NOT_3655(I15814,g11129);
  not NOT_3656(g13251,I15814);
  not NOT_3657(g13255,g10632);
  not NOT_3658(I15821,g11143);
  not NOT_3659(g13258,I15821);
  not NOT_3660(I15824,g1116);
  not NOT_3661(g13259,I15824);
  not NOT_3662(I15831,g10416);
  not NOT_3663(g13267,I15831);
  not NOT_3664(I15834,g11164);
  not NOT_3665(g13271,I15834);
  not NOT_3666(I15837,g1459);
  not NOT_3667(g13272,I15837);
  not NOT_3668(g13278,g10738);
  not NOT_3669(I15843,g11181);
  not NOT_3670(g13279,I15843);
  not NOT_3671(I15846,g11183);
  not NOT_3672(g13280,I15846);
  not NOT_3673(g13297,g10831);
  not NOT_3674(I15862,g11215);
  not NOT_3675(g13298,I15862);
  not NOT_3676(g13301,g10862);
  not NOT_3677(g13302,g12321);
  not NOT_3678(I15869,g11234);
  not NOT_3679(g13303,I15869);
  not NOT_3680(I15872,g11236);
  not NOT_3681(g13304,I15872);
  not NOT_3682(g13305,g11048);
  not NOT_3683(I15878,g11249);
  not NOT_3684(g13311,I15878);
  not NOT_3685(g13312,g11048);
  not NOT_3686(g13314,g10893);
  not NOT_3687(g13322,g10918);
  not NOT_3688(g13323,g11048);
  not NOT_3689(I15893,g10430);
  not NOT_3690(g13329,I15893);
  not NOT_3691(g13334,g11048);
  not NOT_3692(I15906,g10430);
  not NOT_3693(g13350,I15906);
  not NOT_3694(I15915,g10430);
  not NOT_3695(g13394,I15915);
  not NOT_3696(I15918,g12381);
  not NOT_3697(g13409,I15918);
  not NOT_3698(I15921,g12381);
  not NOT_3699(g13410,I15921);
  not NOT_3700(g13412,g11963);
  not NOT_3701(g13413,g11737);
  not NOT_3702(g13414,g11048);
  not NOT_3703(I15929,g10430);
  not NOT_3704(g13416,I15929);
  not NOT_3705(I15932,g12381);
  not NOT_3706(g13431,I15932);
  not NOT_3707(I15937,g11676);
  not NOT_3708(g13437,I15937);
  not NOT_3709(g13458,g11048);
  not NOT_3710(I15942,g12381);
  not NOT_3711(g13460,I15942);
  not NOT_3712(g13463,g10476);
  not NOT_3713(g13474,g11048);
  not NOT_3714(I15954,g12381);
  not NOT_3715(g13477,I15954);
  not NOT_3716(g13483,g11270);
  not NOT_3717(g13484,g10981);
  not NOT_3718(g13485,g10476);
  not NOT_3719(g13494,g11912);
  not NOT_3720(g13504,g11303);
  not NOT_3721(g13505,g10981);
  not NOT_3722(g13506,g10808);
  not NOT_3723(I15981,g11290);
  not NOT_3724(g13510,I15981);
  not NOT_3725(I15987,g12381);
  not NOT_3726(g13514,I15987);
  not NOT_3727(g13521,g11357);
  not NOT_3728(g13522,g10981);
  not NOT_3729(g13530,g12641);
  not NOT_3730(I16010,g11148);
  not NOT_3731(g13545,I16010);
  not NOT_3732(g13555,g12692);
  not NOT_3733(g13565,g11006);
  not NOT_3734(g13569,g10951);
  not NOT_3735(I16024,g11171);
  not NOT_3736(g13574,I16024);
  not NOT_3737(I16028,g12381);
  not NOT_3738(g13583,I16028);
  not NOT_3739(g13584,g12735);
  not NOT_3740(g13593,g10556);
  not NOT_3741(g13594,g11012);
  not NOT_3742(g13595,g10951);
  not NOT_3743(g13596,g10971);
  not NOT_3744(I16040,g10430);
  not NOT_3745(g13605,I16040);
  not NOT_3746(g13620,g10556);
  not NOT_3747(g13621,g10573);
  not NOT_3748(g13624,g10951);
  not NOT_3749(g13625,g10971);
  not NOT_3750(g13626,g11273);
  not NOT_3751(g13637,g10556);
  not NOT_3752(I16057,g10430);
  not NOT_3753(g13638,I16057);
  not NOT_3754(g13655,g10573);
  not NOT_3755(g13663,g10971);
  not NOT_3756(g13664,g11252);
  not NOT_3757(g13665,g11306);
  not NOT_3758(g13675,g10556);
  not NOT_3759(g13679,g10573);
  not NOT_3760(I16077,g10430);
  not NOT_3761(g13680,I16077);
  not NOT_3762(g13706,g11280);
  not NOT_3763(g13707,g11360);
  not NOT_3764(g13715,g10573);
  not NOT_3765(I16090,g10430);
  not NOT_3766(g13716,I16090);
  not NOT_3767(g13729,g10951);
  not NOT_3768(g13736,g11313);
  not NOT_3769(I16102,g10430);
  not NOT_3770(g13745,I16102);
  not NOT_3771(g13763,g10971);
  not NOT_3772(I16117,g10430);
  not NOT_3773(g13782,I16117);
  not NOT_3774(I16120,g11868);
  not NOT_3775(g13793,I16120);
  not NOT_3776(I16135,g10430);
  not NOT_3777(g13809,I16135);
  not NOT_3778(I16150,g10430);
  not NOT_3779(g13835,I16150);
  not NOT_3780(I16160,g11237);
  not NOT_3781(g13856,I16160);
  not NOT_3782(I16163,g11930);
  not NOT_3783(g13857,I16163);
  not NOT_3784(I16168,g3321);
  not NOT_3785(g13865,I16168);
  not NOT_3786(g13868,g11493);
  not NOT_3787(g13869,g10831);
  not NOT_3788(g13876,g11432);
  not NOT_3789(g13877,g11350);
  not NOT_3790(I16181,g3672);
  not NOT_3791(g13881,I16181);
  not NOT_3792(g13885,g10862);
  not NOT_3793(I16193,g3281);
  not NOT_3794(g13895,I16193);
  not NOT_3795(g13901,g11480);
  not NOT_3796(g13902,g11389);
  not NOT_3797(I16201,g4023);
  not NOT_3798(g13906,I16201);
  not NOT_3799(I16217,g3632);
  not NOT_3800(g13926,I16217);
  not NOT_3801(g13932,g11534);
  not NOT_3802(g13933,g11419);
  not NOT_3803(I16231,g10520);
  not NOT_3804(g13943,I16231);
  not NOT_3805(I16246,g3983);
  not NOT_3806(g13966,I16246);
  not NOT_3807(g13975,g11048);
  not NOT_3808(g13976,g11130);
  not NOT_3809(g13995,g11261);
  not NOT_3810(g13999,g11048);
  not NOT_3811(g14004,g11149);
  not NOT_3812(g14029,g11283);
  not NOT_3813(I16289,g12107);
  not NOT_3814(g14031,I16289);
  not NOT_3815(g14032,g11048);
  not NOT_3816(g14034,g11048);
  not NOT_3817(g14063,g11048);
  not NOT_3818(g14065,g11048);
  not NOT_3819(g14095,g11326);
  not NOT_3820(I16328,g878);
  not NOT_3821(g14096,I16328);
  not NOT_3822(I16345,g881);
  not NOT_3823(g14125,I16345);
  not NOT_3824(I16357,g884);
  not NOT_3825(g14147,I16357);
  not NOT_3826(g14149,g12381);
  not NOT_3827(g14150,g12381);
  not NOT_3828(g14166,g11048);
  not NOT_3829(I16371,g887);
  not NOT_3830(g14167,I16371);
  not NOT_3831(g14169,g12381);
  not NOT_3832(g14173,g12076);
  not NOT_3833(g14179,g11048);
  not NOT_3834(g14183,g12381);
  not NOT_3835(g14184,g12381);
  not NOT_3836(g14186,g11346);
  not NOT_3837(I16391,g859);
  not NOT_3838(g14189,I16391);
  not NOT_3839(g14191,g12381);
  not NOT_3840(g14192,g11385);
  not NOT_3841(g14197,g12160);
  not NOT_3842(g14198,g12180);
  not NOT_3843(I16401,g869);
  not NOT_3844(g14201,I16401);
  not NOT_3845(g14203,g12381);
  not NOT_3846(g14204,g12155);
  not NOT_3847(g14205,g12381);
  not NOT_3848(g14208,g11563);
  not NOT_3849(g14209,g11415);
  not NOT_3850(g14215,g12198);
  not NOT_3851(I16417,g875);
  not NOT_3852(g14217,I16417);
  not NOT_3853(g14219,g12381);
  not NOT_3854(g14226,g11618);
  not NOT_3855(g14231,g12246);
  not NOT_3856(g14232,g11083);
  not NOT_3857(g14237,g11666);
  not NOT_3858(g14238,g10823);
  not NOT_3859(g14251,g12308);
  not NOT_3860(I16438,g11165);
  not NOT_3861(g14252,I16438);
  not NOT_3862(g14255,g12381);
  not NOT_3863(g14262,g10838);
  not NOT_3864(g14275,g12358);
  not NOT_3865(I16452,g11182);
  not NOT_3866(g14276,I16452);
  not NOT_3867(I16455,g11845);
  not NOT_3868(g14277,I16455);
  not NOT_3869(I16460,g10430);
  not NOT_3870(g14290,I16460);
  not NOT_3871(g14297,g10869);
  not NOT_3872(I16468,g12760);
  not NOT_3873(g14307,I16468);
  not NOT_3874(I16471,g12367);
  not NOT_3875(g14308,I16471);
  not NOT_3876(I16476,g10430);
  not NOT_3877(g14314,I16476);
  not NOT_3878(I16479,g10430);
  not NOT_3879(g14315,I16479);
  not NOT_3880(g14321,g10874);
  not NOT_3881(I16486,g11204);
  not NOT_3882(g14330,I16486);
  not NOT_3883(I16489,g12793);
  not NOT_3884(g14331,I16489);
  not NOT_3885(I16492,g12430);
  not NOT_3886(g14332,I16492);
  not NOT_3887(I16498,g10430);
  not NOT_3888(g14336,I16498);
  not NOT_3889(I16502,g10430);
  not NOT_3890(g14338,I16502);
  not NOT_3891(g14342,g12163);
  not NOT_3892(g14348,g10887);
  not NOT_3893(g14357,g12181);
  not NOT_3894(I16512,g12811);
  not NOT_3895(g14358,I16512);
  not NOT_3896(I16515,g12477);
  not NOT_3897(g14359,I16515);
  not NOT_3898(I16521,g10430);
  not NOT_3899(g14363,I16521);
  not NOT_3900(I16526,g10430);
  not NOT_3901(g14366,I16526);
  not NOT_3902(g14376,g12126);
  not NOT_3903(g14377,g12201);
  not NOT_3904(I16535,g11235);
  not NOT_3905(g14383,I16535);
  not NOT_3906(I16538,g10417);
  not NOT_3907(g14384,I16538);
  not NOT_3908(I16541,g11929);
  not NOT_3909(g14385,I16541);
  not NOT_3910(I16544,g11931);
  not NOT_3911(g14386,I16544);
  not NOT_3912(I16555,g10430);
  not NOT_3913(g14398,I16555);
  not NOT_3914(g14405,g12170);
  not NOT_3915(g14406,g12249);
  not NOT_3916(I16564,g10429);
  not NOT_3917(g14412,I16564);
  not NOT_3918(I16575,g3298);
  not NOT_3919(g14421,I16575);
  not NOT_3920(I16579,g10981);
  not NOT_3921(g14423,I16579);
  not NOT_3922(g14424,g11136);
  not NOT_3923(g14431,g12208);
  not NOT_3924(g14432,g12311);
  not NOT_3925(I16590,g11966);
  not NOT_3926(g14441,I16590);
  not NOT_3927(I16593,g10498);
  not NOT_3928(g14442,I16593);
  not NOT_3929(I16596,g12640);
  not NOT_3930(g14443,I16596);
  not NOT_3931(I16606,g3649);
  not NOT_3932(g14451,I16606);
  not NOT_3933(I16610,g10981);
  not NOT_3934(g14453,I16610);
  not NOT_3935(I16613,g10430);
  not NOT_3936(g14454,I16613);
  not NOT_3937(g14503,g12256);
  not NOT_3938(g14504,g12361);
  not NOT_3939(I16626,g11986);
  not NOT_3940(g14509,I16626);
  not NOT_3941(I16629,g11987);
  not NOT_3942(g14510,I16629);
  not NOT_3943(I16639,g4000);
  not NOT_3944(g14518,I16639);
  not NOT_3945(g14535,g12318);
  not NOT_3946(I16651,g10542);
  not NOT_3947(g14536,I16651);
  not NOT_3948(g14541,g11405);
  not NOT_3949(I16660,g10981);
  not NOT_3950(g14543,I16660);
  not NOT_3951(I16663,g10981);
  not NOT_3952(g14544,I16663);
  not NOT_3953(g14545,g12768);
  not NOT_3954(g14562,g12036);
  not NOT_3955(I16676,g10588);
  not NOT_3956(g14563,I16676);
  not NOT_3957(I16679,g12039);
  not NOT_3958(g14564,I16679);
  not NOT_3959(I16688,g10981);
  not NOT_3960(g14571,I16688);
  not NOT_3961(I16698,g12077);
  not NOT_3962(g14582,I16698);
  not NOT_3963(g14584,g11048);
  not NOT_3964(I16709,g10430);
  not NOT_3965(g14591,I16709);
  not NOT_3966(I16713,g5331);
  not NOT_3967(g14597,I16713);
  not NOT_3968(I16724,g12108);
  not NOT_3969(g14609,I16724);
  not NOT_3970(I16733,g12026);
  not NOT_3971(g14616,I16733);
  not NOT_3972(g14630,g12402);
  not NOT_3973(g14631,g12239);
  not NOT_3974(I16741,g5677);
  not NOT_3975(g14635,I16741);
  not NOT_3976(I16747,g12729);
  not NOT_3977(g14639,I16747);
  not NOT_3978(I16755,g12377);
  not NOT_3979(g14645,I16755);
  not NOT_3980(I16762,g5290);
  not NOT_3981(g14662,I16762);
  not NOT_3982(g14668,g12450);
  not NOT_3983(g14669,g12301);
  not NOT_3984(I16770,g6023);
  not NOT_3985(g14673,I16770);
  not NOT_3986(I16775,g12183);
  not NOT_3987(g14676,I16775);
  not NOT_3988(I16795,g5637);
  not NOT_3989(g14694,I16795);
  not NOT_3990(g14700,g12512);
  not NOT_3991(g14701,g12351);
  not NOT_3992(I16803,g6369);
  not NOT_3993(g14705,I16803);
  not NOT_3994(g14714,g11405);
  not NOT_3995(I16821,g5983);
  not NOT_3996(g14738,I16821);
  not NOT_3997(g14744,g12578);
  not NOT_3998(g14745,g12423);
  not NOT_3999(I16829,g6715);
  not NOT_4000(g14749,I16829);
  not NOT_4001(g14753,g11317);
  not NOT_4002(I16847,g6329);
  not NOT_4003(g14779,I16847);
  not NOT_4004(g14785,g12629);
  not NOT_4005(g14786,g12471);
  not NOT_4006(I16855,g10473);
  not NOT_4007(g14790,I16855);
  not NOT_4008(I16875,g6675);
  not NOT_4009(g14828,I16875);
  not NOT_4010(g14833,g11405);
  not NOT_4011(I16898,g10615);
  not NOT_4012(g14873,I16898);
  not NOT_4013(I16917,g10582);
  not NOT_4014(g14912,I16917);
  not NOT_4015(I16969,g13943);
  not NOT_4016(g15048,I16969);
  not NOT_4017(I17008,g12857);
  not NOT_4018(g15085,I17008);
  not NOT_4019(I17094,g14331);
  not NOT_4020(g15169,I17094);
  not NOT_4021(I17098,g14336);
  not NOT_4022(g15171,I17098);
  not NOT_4023(I17101,g14338);
  not NOT_4024(g15224,I17101);
  not NOT_4025(I17104,g12932);
  not NOT_4026(g15277,I17104);
  not NOT_4027(g15344,g14851);
  not NOT_4028(I17108,g13782);
  not NOT_4029(g15345,I17108);
  not NOT_4030(I17111,g13809);
  not NOT_4031(g15348,I17111);
  not NOT_4032(I17114,g14358);
  not NOT_4033(g15371,I17114);
  not NOT_4034(I17118,g14363);
  not NOT_4035(g15373,I17118);
  not NOT_4036(I17121,g14366);
  not NOT_4037(g15426,I17121);
  not NOT_4038(g15479,g14895);
  not NOT_4039(I17125,g13809);
  not NOT_4040(g15480,I17125);
  not NOT_4041(I17128,g13835);
  not NOT_4042(g15483,I17128);
  not NOT_4043(I17131,g14384);
  not NOT_4044(g15506,I17131);
  not NOT_4045(I17136,g14398);
  not NOT_4046(g15509,I17136);
  not NOT_4047(g15562,g14943);
  not NOT_4048(I17140,g13835);
  not NOT_4049(g15563,I17140);
  not NOT_4050(I17143,g14412);
  not NOT_4051(g15566,I17143);
  not NOT_4052(g15568,g14984);
  not NOT_4053(I17148,g14442);
  not NOT_4054(g15569,I17148);
  not NOT_4055(g15571,g13211);
  not NOT_4056(I17154,g13605);
  not NOT_4057(g15573,I17154);
  not NOT_4058(I17159,g13350);
  not NOT_4059(g15579,I17159);
  not NOT_4060(g15580,g13242);
  not NOT_4061(I17166,g14536);
  not NOT_4062(g15588,I17166);
  not NOT_4063(I17173,g13716);
  not NOT_4064(g15595,I17173);
  not NOT_4065(g15614,g14914);
  not NOT_4066(I17181,g13745);
  not NOT_4067(g15615,I17181);
  not NOT_4068(I17188,g13782);
  not NOT_4069(g15634,I17188);
  not NOT_4070(g15655,g13202);
  not NOT_4071(I17198,g13809);
  not NOT_4072(g15656,I17198);
  not NOT_4073(I17207,g13835);
  not NOT_4074(g15680,I17207);
  not NOT_4075(g15705,g13217);
  not NOT_4076(I17228,g13350);
  not NOT_4077(g15714,I17228);
  not NOT_4078(g15731,g13326);
  not NOT_4079(I17249,g13605);
  not NOT_4080(g15733,I17249);
  not NOT_4081(g15739,g13284);
  not NOT_4082(g15740,g13342);
  not NOT_4083(g15746,g13121);
  not NOT_4084(g15747,g13307);
  not NOT_4085(g15750,g13291);
  not NOT_4086(g15755,g13134);
  not NOT_4087(g15756,g13315);
  not NOT_4088(I17276,g13605);
  not NOT_4089(g15758,I17276);
  not NOT_4090(g15799,g13110);
  not NOT_4091(I17302,g14044);
  not NOT_4092(g15806,I17302);
  not NOT_4093(g15811,g13125);
  not NOT_4094(I17314,g14078);
  not NOT_4095(g15816,I17314);
  not NOT_4096(I17324,g14119);
  not NOT_4097(g15824,I17324);
  not NOT_4098(g15830,g13432);
  not NOT_4099(g15831,g13385);
  not NOT_4100(g15842,g13469);
  not NOT_4101(I17355,g14591);
  not NOT_4102(g15862,I17355);
  not NOT_4103(I17374,g13638);
  not NOT_4104(g15885,I17374);
  not NOT_4105(I17392,g13680);
  not NOT_4106(g15915,I17392);
  not NOT_4107(I17395,g12952);
  not NOT_4108(g15932,I17395);
  not NOT_4109(I17401,g13394);
  not NOT_4110(g15938,I17401);
  not NOT_4111(I17416,g13806);
  not NOT_4112(g15969,I17416);
  not NOT_4113(I17420,g13394);
  not NOT_4114(g15979,I17420);
  not NOT_4115(I17425,g13416);
  not NOT_4116(g16000,I17425);
  not NOT_4117(g16030,g13570);
  not NOT_4118(I17436,g13416);
  not NOT_4119(g16031,I17436);
  not NOT_4120(I17442,g13638);
  not NOT_4121(g16053,I17442);
  not NOT_4122(g16075,g13597);
  not NOT_4123(I17456,g13680);
  not NOT_4124(g16077,I17456);
  not NOT_4125(g16096,g13530);
  not NOT_4126(g16099,g13437);
  not NOT_4127(I17471,g13394);
  not NOT_4128(g16100,I17471);
  not NOT_4129(g16123,g13530);
  not NOT_4130(g16124,g13555);
  not NOT_4131(g16127,g13437);
  not NOT_4132(I17488,g13394);
  not NOT_4133(g16129,I17488);
  not NOT_4134(I17491,g13416);
  not NOT_4135(g16136,I17491);
  not NOT_4136(g16158,g13555);
  not NOT_4137(g16159,g13584);
  not NOT_4138(g16162,g13437);
  not NOT_4139(I17507,g13416);
  not NOT_4140(g16164,I17507);
  not NOT_4141(g16171,g13530);
  not NOT_4142(g16172,g13584);
  not NOT_4143(g16180,g13437);
  not NOT_4144(g16182,g13846);
  not NOT_4145(g16186,g13555);
  not NOT_4146(g16195,g13437);
  not NOT_4147(g16197,g13861);
  not NOT_4148(g16200,g13584);
  not NOT_4149(g16206,g13437);
  not NOT_4150(g16214,g13437);
  not NOT_4151(I17557,g14510);
  not NOT_4152(g16216,I17557);
  not NOT_4153(g16223,g13437);
  not NOT_4154(I17569,g14564);
  not NOT_4155(g16228,I17569);
  not NOT_4156(g16235,g13437);
  not NOT_4157(I17590,g14591);
  not NOT_4158(g16249,I17590);
  not NOT_4159(g16280,g13330);
  not NOT_4160(I17609,g13510);
  not NOT_4161(g16284,I17609);
  not NOT_4162(I17612,g13250);
  not NOT_4163(g16285,I17612);
  not NOT_4164(I17615,g13251);
  not NOT_4165(g16286,I17615);
  not NOT_4166(g16289,g13223);
  not NOT_4167(g16290,g13260);
  not NOT_4168(I17626,g14582);
  not NOT_4169(g16300,I17626);
  not NOT_4170(g16305,g13346);
  not NOT_4171(I17633,g13258);
  not NOT_4172(g16307,I17633);
  not NOT_4173(I17636,g14252);
  not NOT_4174(g16308,I17636);
  not NOT_4175(I17639,g13350);
  not NOT_4176(g16309,I17639);
  not NOT_4177(g16310,g13223);
  not NOT_4178(g16311,g13273);
  not NOT_4179(g16320,g14454);
  not NOT_4180(I17650,g13271);
  not NOT_4181(g16322,I17650);
  not NOT_4182(I17653,g14276);
  not NOT_4183(g16323,I17653);
  not NOT_4184(g16325,g13223);
  not NOT_4185(I17658,g13394);
  not NOT_4186(g16326,I17658);
  not NOT_4187(I17661,g13329);
  not NOT_4188(g16349,I17661);
  not NOT_4189(g16423,g14066);
  not NOT_4190(I17668,g13279);
  not NOT_4191(g16428,I17668);
  not NOT_4192(I17671,g13280);
  not NOT_4193(g16429,I17671);
  not NOT_4194(I17675,g13394);
  not NOT_4195(g16431,I17675);
  not NOT_4196(I17679,g13416);
  not NOT_4197(g16449,I17679);
  not NOT_4198(g16472,g14098);
  not NOT_4199(g16473,g13977);
  not NOT_4200(g16475,g14107);
  not NOT_4201(g16482,g13464);
  not NOT_4202(I17695,g14330);
  not NOT_4203(g16487,I17695);
  not NOT_4204(I17699,g13416);
  not NOT_4205(g16489,I17699);
  not NOT_4206(I17704,g13144);
  not NOT_4207(g16508,I17704);
  not NOT_4208(g16509,g13873);
  not NOT_4209(g16510,g14008);
  not NOT_4210(g16511,g14130);
  not NOT_4211(g16512,g14015);
  not NOT_4212(g16514,g14139);
  not NOT_4213(g16515,g13486);
  not NOT_4214(g16521,g13543);
  not NOT_4215(g16522,g13889);
  not NOT_4216(g16523,g14041);
  not NOT_4217(I17723,g13177);
  not NOT_4218(g16525,I17723);
  not NOT_4219(g16526,g13898);
  not NOT_4220(g16527,g14048);
  not NOT_4221(g16528,g14154);
  not NOT_4222(g16529,g14055);
  not NOT_4223(g16530,g14454);
  not NOT_4224(I17733,g14844);
  not NOT_4225(g16533,I17733);
  not NOT_4226(I17744,g14912);
  not NOT_4227(g16540,I17744);
  not NOT_4228(I17747,g13298);
  not NOT_4229(g16577,I17747);
  not NOT_4230(I17750,g14383);
  not NOT_4231(g16578,I17750);
  not NOT_4232(g16579,g13267);
  not NOT_4233(I17754,g13494);
  not NOT_4234(g16580,I17754);
  not NOT_4235(g16582,g13915);
  not NOT_4236(g16583,g14069);
  not NOT_4237(g16584,g13920);
  not NOT_4238(g16585,g14075);
  not NOT_4239(I17763,g13191);
  not NOT_4240(g16587,I17763);
  not NOT_4241(g16588,g13929);
  not NOT_4242(g16589,g14082);
  not NOT_4243(I17772,g14888);
  not NOT_4244(g16594,I17772);
  not NOT_4245(I17780,g13303);
  not NOT_4246(g16600,I17780);
  not NOT_4247(I17783,g13304);
  not NOT_4248(g16601,I17783);
  not NOT_4249(g16602,g14101);
  not NOT_4250(I17787,g3267);
  not NOT_4251(g16603,I17787);
  not NOT_4252(g16605,g13955);
  not NOT_4253(g16606,g14110);
  not NOT_4254(g16607,g13960);
  not NOT_4255(g16608,g14116);
  not NOT_4256(g16609,g14454);
  not NOT_4257(I17801,g14936);
  not NOT_4258(g16615,I17801);
  not NOT_4259(I17808,g13311);
  not NOT_4260(g16620,I17808);
  not NOT_4261(g16622,g14104);
  not NOT_4262(g16623,g14127);
  not NOT_4263(I17814,g3274);
  not NOT_4264(g16624,I17814);
  not NOT_4265(g16626,g14133);
  not NOT_4266(I17819,g3618);
  not NOT_4267(g16627,I17819);
  not NOT_4268(g16629,g13990);
  not NOT_4269(g16630,g14142);
  not NOT_4270(g16631,g14454);
  not NOT_4271(g16632,g14454);
  not NOT_4272(I17834,g14977);
  not NOT_4273(g16640,I17834);
  not NOT_4274(I17839,g13412);
  not NOT_4275(g16643,I17839);
  not NOT_4276(I17842,g13051);
  not NOT_4277(g16644,I17842);
  not NOT_4278(g16645,g13756);
  not NOT_4279(g16651,g14005);
  not NOT_4280(g16652,g13892);
  not NOT_4281(g16654,g14136);
  not NOT_4282(g16655,g14151);
  not NOT_4283(I17852,g3625);
  not NOT_4284(g16656,I17852);
  not NOT_4285(g16658,g14157);
  not NOT_4286(I17857,g3969);
  not NOT_4287(g16659,I17857);
  not NOT_4288(g16661,g14454);
  not NOT_4289(I17873,g15017);
  not NOT_4290(g16675,I17873);
  not NOT_4291(I17876,g13070);
  not NOT_4292(g16676,I17876);
  not NOT_4293(I17879,g14386);
  not NOT_4294(g16677,I17879);
  not NOT_4295(g16680,g13223);
  not NOT_4296(g16684,g14223);
  not NOT_4297(g16685,g14038);
  not NOT_4298(I17892,g3325);
  not NOT_4299(g16686,I17892);
  not NOT_4300(g16688,g14045);
  not NOT_4301(g16689,g13923);
  not NOT_4302(g16691,g14160);
  not NOT_4303(g16692,g14170);
  not NOT_4304(I17901,g3976);
  not NOT_4305(g16693,I17901);
  not NOT_4306(g16695,g14454);
  not NOT_4307(I17916,g13087);
  not NOT_4308(g16708,I17916);
  not NOT_4309(I17919,g14609);
  not NOT_4310(g16709,I17919);
  not NOT_4311(g16712,g13223);
  not NOT_4312(g16716,g13948);
  not NOT_4313(g16717,g13951);
  not NOT_4314(I17932,g3310);
  not NOT_4315(g16718,I17932);
  not NOT_4316(g16720,g14234);
  not NOT_4317(g16721,g14072);
  not NOT_4318(I17938,g3676);
  not NOT_4319(g16722,I17938);
  not NOT_4320(g16724,g14079);
  not NOT_4321(g16725,g13963);
  not NOT_4322(g16726,g14454);
  not NOT_4323(g16727,g14454);
  not NOT_4324(I17956,g14562);
  not NOT_4325(g16738,I17956);
  not NOT_4326(g16739,g13223);
  not NOT_4327(g16740,g13980);
  not NOT_4328(g16742,g13983);
  not NOT_4329(g16743,g13986);
  not NOT_4330(I17964,g3661);
  not NOT_4331(g16744,I17964);
  not NOT_4332(g16746,g14258);
  not NOT_4333(g16747,g14113);
  not NOT_4334(I17970,g4027);
  not NOT_4335(g16748,I17970);
  not NOT_4336(g16750,g14454);
  not NOT_4337(I17976,g13638);
  not NOT_4338(g16752,I17976);
  not NOT_4339(I17989,g14173);
  not NOT_4340(g16767,I17989);
  not NOT_4341(g16768,g13223);
  not NOT_4342(g16769,g13530);
  not NOT_4343(g16771,g14018);
  not NOT_4344(g16773,g14021);
  not NOT_4345(g16774,g14024);
  not NOT_4346(I17999,g4012);
  not NOT_4347(g16775,I17999);
  not NOT_4348(I18003,g13638);
  not NOT_4349(g16777,I18003);
  not NOT_4350(I18006,g13638);
  not NOT_4351(g16782,I18006);
  not NOT_4352(I18009,g13680);
  not NOT_4353(g16795,I18009);
  not NOT_4354(g16809,g14387);
  not NOT_4355(g16812,g13555);
  not NOT_4356(g16814,g14058);
  not NOT_4357(I18028,g13638);
  not NOT_4358(g16816,I18028);
  not NOT_4359(I18031,g13680);
  not NOT_4360(g16821,I18031);
  not NOT_4361(I18034,g13680);
  not NOT_4362(g16826,I18034);
  not NOT_4363(g16853,g13584);
  not NOT_4364(I18048,g13638);
  not NOT_4365(g16856,I18048);
  not NOT_4366(I18051,g13680);
  not NOT_4367(g16861,I18051);
  not NOT_4368(I18060,g14198);
  not NOT_4369(g16872,I18060);
  not NOT_4370(I18063,g14357);
  not NOT_4371(g16873,I18063);
  not NOT_4372(I18066,g3317);
  not NOT_4373(g16874,I18066);
  not NOT_4374(I18071,g13680);
  not NOT_4375(g16877,I18071);
  not NOT_4376(I18078,g13350);
  not NOT_4377(g16886,I18078);
  not NOT_4378(I18083,g13394);
  not NOT_4379(g16897,I18083);
  not NOT_4380(I18086,g13856);
  not NOT_4381(g16920,I18086);
  not NOT_4382(I18089,g13144);
  not NOT_4383(g16923,I18089);
  not NOT_4384(I18092,g3668);
  not NOT_4385(g16924,I18092);
  not NOT_4386(I18101,g13416);
  not NOT_4387(g16931,I18101);
  not NOT_4388(I18104,g13177);
  not NOT_4389(g16954,I18104);
  not NOT_4390(I18107,g4019);
  not NOT_4391(g16955,I18107);
  not NOT_4392(g16958,g14238);
  not NOT_4393(I18114,g14509);
  not NOT_4394(g16960,I18114);
  not NOT_4395(I18117,g13302);
  not NOT_4396(g16963,I18117);
  not NOT_4397(I18120,g13350);
  not NOT_4398(g16964,I18120);
  not NOT_4399(g16966,g14291);
  not NOT_4400(I18125,g13191);
  not NOT_4401(g16967,I18125);
  not NOT_4402(g16968,g14238);
  not NOT_4403(g16969,g14262);
  not NOT_4404(I18131,g13350);
  not NOT_4405(g16971,I18131);
  not NOT_4406(I18135,g13144);
  not NOT_4407(g16987,I18135);
  not NOT_4408(I18138,g14277);
  not NOT_4409(g17010,I18138);
  not NOT_4410(g17013,g14262);
  not NOT_4411(g17014,g14297);
  not NOT_4412(I18143,g13350);
  not NOT_4413(g17015,I18143);
  not NOT_4414(g17056,g13437);
  not NOT_4415(I18148,g13526);
  not NOT_4416(g17058,I18148);
  not NOT_4417(I18151,g13144);
  not NOT_4418(g17059,I18151);
  not NOT_4419(I18154,g13177);
  not NOT_4420(g17062,I18154);
  not NOT_4421(g17085,g14238);
  not NOT_4422(g17086,g14297);
  not NOT_4423(g17087,g14321);
  not NOT_4424(I18160,g14441);
  not NOT_4425(g17088,I18160);
  not NOT_4426(g17092,g14011);
  not NOT_4427(I18165,g13177);
  not NOT_4428(g17093,I18165);
  not NOT_4429(I18168,g13191);
  not NOT_4430(g17096,I18168);
  not NOT_4431(g17120,g14262);
  not NOT_4432(g17121,g14321);
  not NOT_4433(g17122,g14348);
  not NOT_4434(g17124,g14051);
  not NOT_4435(I18177,g13191);
  not NOT_4436(g17125,I18177);
  not NOT_4437(I18180,g13605);
  not NOT_4438(g17128,I18180);
  not NOT_4439(g17135,g14297);
  not NOT_4440(g17136,g14348);
  not NOT_4441(I18191,g14385);
  not NOT_4442(g17141,I18191);
  not NOT_4443(g17144,g14085);
  not NOT_4444(g17147,g14321);
  not NOT_4445(g17154,g14348);
  not NOT_4446(I18205,g14563);
  not NOT_4447(g17155,I18205);
  not NOT_4448(g17157,g13350);
  not NOT_4449(I18214,g12918);
  not NOT_4450(g17178,I18214);
  not NOT_4451(I18221,g13605);
  not NOT_4452(g17183,I18221);
  not NOT_4453(I18224,g13793);
  not NOT_4454(g17188,I18224);
  not NOT_4455(g17189,g14708);
  not NOT_4456(I18233,g14639);
  not NOT_4457(g17197,I18233);
  not NOT_4458(I18238,g13144);
  not NOT_4459(g17200,I18238);
  not NOT_4460(g17216,g14454);
  not NOT_4461(I18245,g14676);
  not NOT_4462(g17221,I18245);
  not NOT_4463(I18248,g12938);
  not NOT_4464(g17224,I18248);
  not NOT_4465(I18252,g13177);
  not NOT_4466(g17226,I18252);
  not NOT_4467(g17242,g14454);
  not NOT_4468(I18259,g12946);
  not NOT_4469(g17247,I18259);
  not NOT_4470(I18262,g13857);
  not NOT_4471(g17248,I18262);
  not NOT_4472(I18265,g13350);
  not NOT_4473(g17249,I18265);
  not NOT_4474(I18270,g13191);
  not NOT_4475(g17271,I18270);
  not NOT_4476(I18276,g1075);
  not NOT_4477(g17291,I18276);
  not NOT_4478(I18280,g12951);
  not NOT_4479(g17296,I18280);
  not NOT_4480(g17301,g14454);
  not NOT_4481(I18285,g13638);
  not NOT_4482(g17302,I18285);
  not NOT_4483(g17308,g14876);
  not NOT_4484(I18293,g1079);
  not NOT_4485(g17316,I18293);
  not NOT_4486(I18297,g1418);
  not NOT_4487(g17320,I18297);
  not NOT_4488(I18301,g12976);
  not NOT_4489(g17324,I18301);
  not NOT_4490(I18304,g14790);
  not NOT_4491(g17325,I18304);
  not NOT_4492(I18307,g12977);
  not NOT_4493(g17326,I18307);
  not NOT_4494(I18310,g12978);
  not NOT_4495(g17327,I18310);
  not NOT_4496(I18313,g13350);
  not NOT_4497(g17328,I18313);
  not NOT_4498(g17366,g14454);
  not NOT_4499(I18320,g13605);
  not NOT_4500(g17367,I18320);
  not NOT_4501(I18323,g13680);
  not NOT_4502(g17384,I18323);
  not NOT_4503(g17389,g14915);
  not NOT_4504(g17390,g14755);
  not NOT_4505(g17392,g14924);
  not NOT_4506(I18333,g1083);
  not NOT_4507(g17400,I18333);
  not NOT_4508(I18337,g1422);
  not NOT_4509(g17404,I18337);
  not NOT_4510(I18341,g14308);
  not NOT_4511(g17408,I18341);
  not NOT_4512(I18344,g13003);
  not NOT_4513(g17409,I18344);
  not NOT_4514(g17410,g12955);
  not NOT_4515(g17411,g14454);
  not NOT_4516(I18350,g13716);
  not NOT_4517(g17413,I18350);
  not NOT_4518(g17414,g14627);
  not NOT_4519(g17415,g14797);
  not NOT_4520(g17416,g14956);
  not NOT_4521(g17417,g14804);
  not NOT_4522(g17419,g14965);
  not NOT_4523(I18360,g1426);
  not NOT_4524(g17423,I18360);
  not NOT_4525(I18364,g13009);
  not NOT_4526(g17427,I18364);
  not NOT_4527(I18367,g13010);
  not NOT_4528(g17428,I18367);
  not NOT_4529(I18370,g14873);
  not NOT_4530(g17429,I18370);
  not NOT_4531(I18373,g13011);
  not NOT_4532(g17430,I18373);
  not NOT_4533(I18376,g14332);
  not NOT_4534(g17431,I18376);
  not NOT_4535(I18379,g13012);
  not NOT_4536(g17432,I18379);
  not NOT_4537(I18382,g13350);
  not NOT_4538(g17433,I18382);
  not NOT_4539(g17465,g12955);
  not NOT_4540(g17466,g12983);
  not NOT_4541(g17467,g14339);
  not NOT_4542(g17470,g14454);
  not NOT_4543(g17471,g14454);
  not NOT_4544(g17472,g14656);
  not NOT_4545(g17473,g14841);
  not NOT_4546(I18398,g13745);
  not NOT_4547(g17475,I18398);
  not NOT_4548(g17476,g14665);
  not NOT_4549(g17477,g14848);
  not NOT_4550(g17478,g14996);
  not NOT_4551(g17479,g14855);
  not NOT_4552(g17481,g15005);
  not NOT_4553(I18408,g13017);
  not NOT_4554(g17485,I18408);
  not NOT_4555(I18411,g13018);
  not NOT_4556(g17486,I18411);
  not NOT_4557(I18414,g14359);
  not NOT_4558(g17487,I18414);
  not NOT_4559(g17489,g12955);
  not NOT_4560(g17491,g12983);
  not NOT_4561(g17494,g14339);
  not NOT_4562(g17496,g14683);
  not NOT_4563(g17497,g14879);
  not NOT_4564(g17498,g14688);
  not NOT_4565(g17499,g14885);
  not NOT_4566(I18434,g13782);
  not NOT_4567(g17501,I18434);
  not NOT_4568(g17502,g14697);
  not NOT_4569(g17503,g14892);
  not NOT_4570(g17504,g15021);
  not NOT_4571(g17505,g14899);
  not NOT_4572(g17507,g15030);
  not NOT_4573(I18443,g13027);
  not NOT_4574(g17508,I18443);
  not NOT_4575(I18446,g13028);
  not NOT_4576(g17509,I18446);
  not NOT_4577(g17512,g12983);
  not NOT_4578(g17518,g14918);
  not NOT_4579(I18460,g5276);
  not NOT_4580(g17519,I18460);
  not NOT_4581(g17521,g14727);
  not NOT_4582(g17522,g14927);
  not NOT_4583(g17523,g14732);
  not NOT_4584(g17524,g14933);
  not NOT_4585(I18469,g13809);
  not NOT_4586(g17526,I18469);
  not NOT_4587(g17527,g14741);
  not NOT_4588(g17528,g14940);
  not NOT_4589(g17529,g15039);
  not NOT_4590(g17530,g14947);
  not NOT_4591(I18476,g14031);
  not NOT_4592(g17531,I18476);
  not NOT_4593(I18479,g13041);
  not NOT_4594(g17532,I18479);
  not NOT_4595(I18482,g13350);
  not NOT_4596(g17533,I18482);
  not NOT_4597(g17573,g12911);
  not NOT_4598(g17575,g14921);
  not NOT_4599(g17576,g14953);
  not NOT_4600(I18504,g5283);
  not NOT_4601(g17577,I18504);
  not NOT_4602(g17579,g14959);
  not NOT_4603(I18509,g5623);
  not NOT_4604(g17580,I18509);
  not NOT_4605(g17582,g14768);
  not NOT_4606(g17583,g14968);
  not NOT_4607(g17584,g14773);
  not NOT_4608(g17585,g14974);
  not NOT_4609(I18518,g13835);
  not NOT_4610(g17587,I18518);
  not NOT_4611(g17588,g14782);
  not NOT_4612(g17589,g14981);
  not NOT_4613(I18523,g14443);
  not NOT_4614(g17590,I18523);
  not NOT_4615(I18526,g13055);
  not NOT_4616(g17591,I18526);
  not NOT_4617(g17599,g14794);
  not NOT_4618(g17600,g14659);
  not NOT_4619(g17602,g14962);
  not NOT_4620(g17603,g14993);
  not NOT_4621(I18555,g5630);
  not NOT_4622(g17604,I18555);
  not NOT_4623(g17606,g14999);
  not NOT_4624(I18560,g5969);
  not NOT_4625(g17607,I18560);
  not NOT_4626(g17609,g14817);
  not NOT_4627(g17610,g15008);
  not NOT_4628(g17611,g14822);
  not NOT_4629(g17612,g15014);
  not NOT_4630(I18571,g13074);
  not NOT_4631(g17614,I18571);
  not NOT_4632(I18574,g13075);
  not NOT_4633(g17615,I18574);
  not NOT_4634(g17616,g14309);
  not NOT_4635(g17637,g12933);
  not NOT_4636(g17638,g14838);
  not NOT_4637(I18600,g5335);
  not NOT_4638(g17639,I18600);
  not NOT_4639(g17641,g14845);
  not NOT_4640(g17642,g14691);
  not NOT_4641(g17644,g15002);
  not NOT_4642(g17645,g15018);
  not NOT_4643(I18609,g5976);
  not NOT_4644(g17646,I18609);
  not NOT_4645(g17648,g15024);
  not NOT_4646(I18614,g6315);
  not NOT_4647(g17649,I18614);
  not NOT_4648(g17651,g14868);
  not NOT_4649(g17652,g15033);
  not NOT_4650(g17672,g14720);
  not NOT_4651(g17673,g14723);
  not NOT_4652(I18647,g5320);
  not NOT_4653(g17674,I18647);
  not NOT_4654(g17676,g12941);
  not NOT_4655(g17677,g14882);
  not NOT_4656(I18653,g5681);
  not NOT_4657(g17678,I18653);
  not NOT_4658(g17680,g14889);
  not NOT_4659(g17681,g14735);
  not NOT_4660(g17683,g15027);
  not NOT_4661(g17684,g15036);
  not NOT_4662(I18662,g6322);
  not NOT_4663(g17685,I18662);
  not NOT_4664(g17687,g15042);
  not NOT_4665(I18667,g6661);
  not NOT_4666(g17688,I18667);
  not NOT_4667(I18674,g13101);
  not NOT_4668(g17691,I18674);
  not NOT_4669(g17707,g14758);
  not NOT_4670(g17709,g14761);
  not NOT_4671(g17710,g14764);
  not NOT_4672(I18694,g5666);
  not NOT_4673(g17711,I18694);
  not NOT_4674(g17713,g12947);
  not NOT_4675(g17714,g14930);
  not NOT_4676(I18700,g6027);
  not NOT_4677(g17715,I18700);
  not NOT_4678(g17717,g14937);
  not NOT_4679(g17718,g14776);
  not NOT_4680(g17720,g15045);
  not NOT_4681(g17721,g12915);
  not NOT_4682(I18709,g6668);
  not NOT_4683(g17722,I18709);
  not NOT_4684(g17733,g14238);
  not NOT_4685(g17735,g14807);
  not NOT_4686(g17737,g14810);
  not NOT_4687(g17738,g14813);
  not NOT_4688(I18728,g6012);
  not NOT_4689(g17739,I18728);
  not NOT_4690(g17741,g12972);
  not NOT_4691(g17742,g14971);
  not NOT_4692(I18734,g6373);
  not NOT_4693(g17743,I18734);
  not NOT_4694(g17745,g14978);
  not NOT_4695(g17746,g14825);
  not NOT_4696(g17754,g14262);
  not NOT_4697(g17756,g14858);
  not NOT_4698(g17758,g14861);
  not NOT_4699(g17759,g14864);
  not NOT_4700(I18752,g6358);
  not NOT_4701(g17760,I18752);
  not NOT_4702(g17762,g13000);
  not NOT_4703(g17763,g15011);
  not NOT_4704(I18758,g6719);
  not NOT_4705(g17764,I18758);
  not NOT_4706(g17772,g14297);
  not NOT_4707(g17774,g14902);
  not NOT_4708(g17776,g14905);
  not NOT_4709(g17777,g14908);
  not NOT_4710(I18778,g6704);
  not NOT_4711(g17778,I18778);
  not NOT_4712(I18788,g13138);
  not NOT_4713(g17782,I18788);
  not NOT_4714(I18795,g5327);
  not NOT_4715(g17787,I18795);
  not NOT_4716(g17789,g14321);
  not NOT_4717(g17791,g14950);
  not NOT_4718(g17794,g13350);
  not NOT_4719(g17811,g12925);
  not NOT_4720(I18810,g13716);
  not NOT_4721(g17812,I18810);
  not NOT_4722(I18813,g5673);
  not NOT_4723(g17813,I18813);
  not NOT_4724(g17815,g14348);
  not NOT_4725(I18822,g13745);
  not NOT_4726(g17818,I18822);
  not NOT_4727(I18825,g6019);
  not NOT_4728(g17819,I18825);
  not NOT_4729(I18829,g13350);
  not NOT_4730(g17821,I18829);
  not NOT_4731(I18832,g13782);
  not NOT_4732(g17844,I18832);
  not NOT_4733(I18835,g6365);
  not NOT_4734(g17845,I18835);
  not NOT_4735(I18839,g13716);
  not NOT_4736(g17847,I18839);
  not NOT_4737(I18842,g13809);
  not NOT_4738(g17870,I18842);
  not NOT_4739(I18845,g6711);
  not NOT_4740(g17871,I18845);
  not NOT_4741(I18849,g14290);
  not NOT_4742(g17873,I18849);
  not NOT_4743(I18852,g13716);
  not NOT_4744(g17926,I18852);
  not NOT_4745(I18855,g13745);
  not NOT_4746(g17929,I18855);
  not NOT_4747(I18858,g13835);
  not NOT_4748(g17952,I18858);
  not NOT_4749(I18861,g14307);
  not NOT_4750(g17953,I18861);
  not NOT_4751(I18865,g14314);
  not NOT_4752(g17955,I18865);
  not NOT_4753(I18868,g14315);
  not NOT_4754(g18008,I18868);
  not NOT_4755(g18061,g14800);
  not NOT_4756(I18872,g13745);
  not NOT_4757(g18062,I18872);
  not NOT_4758(I18875,g13782);
  not NOT_4759(g18065,I18875);
  not NOT_4760(g18088,g13267);
  not NOT_4761(I18879,g13267);
  not NOT_4762(g18091,I18879);
  not NOT_4763(I18882,g16580);
  not NOT_4764(g18092,I18882);
  not NOT_4765(I18885,g16643);
  not NOT_4766(g18093,I18885);
  not NOT_4767(I18888,g16644);
  not NOT_4768(g18094,I18888);
  not NOT_4769(I18891,g16676);
  not NOT_4770(g18095,I18891);
  not NOT_4771(I18894,g16708);
  not NOT_4772(g18096,I18894);
  not NOT_4773(I18897,g16738);
  not NOT_4774(g18097,I18897);
  not NOT_4775(I18900,g16767);
  not NOT_4776(g18098,I18900);
  not NOT_4777(I18903,g16872);
  not NOT_4778(g18099,I18903);
  not NOT_4779(I18906,g16963);
  not NOT_4780(g18100,I18906);
  not NOT_4781(I18909,g16873);
  not NOT_4782(g18101,I18909);
  not NOT_4783(I18912,g15050);
  not NOT_4784(g18102,I18912);
  not NOT_4785(I19012,g15060);
  not NOT_4786(g18200,I19012);
  not NOT_4787(I19235,g15078);
  not NOT_4788(g18421,I19235);
  not NOT_4789(I19238,g15079);
  not NOT_4790(g18422,I19238);
  not NOT_4791(I19345,g15083);
  not NOT_4792(g18527,I19345);
  not NOT_4793(I19348,g15084);
  not NOT_4794(g18528,I19348);
  not NOT_4795(I19384,g15085);
  not NOT_4796(g18562,I19384);
  not NOT_4797(I19484,g15122);
  not NOT_4798(g18660,I19484);
  not NOT_4799(I19487,g15125);
  not NOT_4800(g18661,I19487);
  not NOT_4801(g18827,g16000);
  not NOT_4802(g18828,g17955);
  not NOT_4803(g18829,g15171);
  not NOT_4804(g18830,g18008);
  not NOT_4805(g18831,g15224);
  not NOT_4806(g18832,g15634);
  not NOT_4807(I19661,g17587);
  not NOT_4808(g18833,I19661);
  not NOT_4809(g18874,g15938);
  not NOT_4810(g18875,g15171);
  not NOT_4811(g18876,g15373);
  not NOT_4812(g18877,g15224);
  not NOT_4813(g18878,g15426);
  not NOT_4814(g18880,g15656);
  not NOT_4815(I19671,g15932);
  not NOT_4816(g18881,I19671);
  not NOT_4817(I19674,g15932);
  not NOT_4818(g18882,I19674);
  not NOT_4819(g18883,g15938);
  not NOT_4820(g18884,g15938);
  not NOT_4821(g18885,g15979);
  not NOT_4822(g18886,g16000);
  not NOT_4823(g18887,g15373);
  not NOT_4824(g18888,g15426);
  not NOT_4825(g18889,g15509);
  not NOT_4826(g18891,g16053);
  not NOT_4827(g18892,g15680);
  not NOT_4828(g18894,g16000);
  not NOT_4829(g18895,g16000);
  not NOT_4830(g18896,g16031);
  not NOT_4831(g18897,g15509);
  not NOT_4832(g18898,g15566);
  not NOT_4833(g18903,g15758);
  not NOT_4834(g18904,g16053);
  not NOT_4835(g18905,g16077);
  not NOT_4836(g18907,g15979);
  not NOT_4837(g18908,g16100);
  not NOT_4838(g18911,g15169);
  not NOT_4839(g18916,g16053);
  not NOT_4840(g18917,g16077);
  not NOT_4841(I19704,g17653);
  not NOT_4842(g18918,I19704);
  not NOT_4843(I19707,g17590);
  not NOT_4844(g18926,I19707);
  not NOT_4845(g18929,g16100);
  not NOT_4846(g18930,g15789);
  not NOT_4847(g18931,g16031);
  not NOT_4848(g18932,g16136);
  not NOT_4849(g18938,g16053);
  not NOT_4850(g18939,g16077);
  not NOT_4851(I19719,g17431);
  not NOT_4852(g18940,I19719);
  not NOT_4853(g18944,g15938);
  not NOT_4854(g18945,g16100);
  not NOT_4855(g18946,g16100);
  not NOT_4856(g18947,g16136);
  not NOT_4857(g18948,g15800);
  not NOT_4858(g18952,g16053);
  not NOT_4859(g18953,g16077);
  not NOT_4860(g18954,g17427);
  not NOT_4861(I19734,g17725);
  not NOT_4862(g18957,I19734);
  not NOT_4863(g18975,g15938);
  not NOT_4864(g18976,g16100);
  not NOT_4865(g18977,g16100);
  not NOT_4866(g18978,g16000);
  not NOT_4867(g18979,g16136);
  not NOT_4868(g18980,g16136);
  not NOT_4869(g18983,g16077);
  not NOT_4870(g18984,g17486);
  not NOT_4871(g18988,g15979);
  not NOT_4872(g18989,g16000);
  not NOT_4873(g18990,g16136);
  not NOT_4874(g18991,g16136);
  not NOT_4875(I19756,g17812);
  not NOT_4876(g18997,I19756);
  not NOT_4877(I19759,g17767);
  not NOT_4878(g19050,I19759);
  not NOT_4879(I19762,g15732);
  not NOT_4880(g19061,I19762);
  not NOT_4881(g19067,g15979);
  not NOT_4882(g19068,g16031);
  not NOT_4883(g19071,g15591);
  not NOT_4884(I19772,g17818);
  not NOT_4885(g19074,I19772);
  not NOT_4886(I19775,g17780);
  not NOT_4887(g19127,I19775);
  not NOT_4888(I19778,g17781);
  not NOT_4889(g19128,I19778);
  not NOT_4890(g19144,g16031);
  not NOT_4891(g19146,g15574);
  not NOT_4892(I19786,g17844);
  not NOT_4893(g19147,I19786);
  not NOT_4894(I19789,g17793);
  not NOT_4895(g19200,I19789);
  not NOT_4896(g19208,g17367);
  not NOT_4897(I19796,g17870);
  not NOT_4898(g19210,I19796);
  not NOT_4899(I19799,g17817);
  not NOT_4900(g19263,I19799);
  not NOT_4901(I19802,g15727);
  not NOT_4902(g19264,I19802);
  not NOT_4903(g19273,g16100);
  not NOT_4904(g19276,g17367);
  not NOT_4905(I19813,g17952);
  not NOT_4906(g19277,I19813);
  not NOT_4907(g19330,g17326);
  not NOT_4908(I19818,g1056);
  not NOT_4909(g19334,I19818);
  not NOT_4910(g19343,g16136);
  not NOT_4911(g19345,g17591);
  not NOT_4912(g19351,g17367);
  not NOT_4913(g19352,g15758);
  not NOT_4914(I19831,g16533);
  not NOT_4915(g19353,I19831);
  not NOT_4916(g19355,g16027);
  not NOT_4917(I19837,g1399);
  not NOT_4918(g19357,I19837);
  not NOT_4919(g19360,g16249);
  not NOT_4920(I19843,g16594);
  not NOT_4921(g19361,I19843);
  not NOT_4922(g19362,g16072);
  not NOT_4923(g19364,g15825);
  not NOT_4924(g19365,g16249);
  not NOT_4925(g19366,g15885);
  not NOT_4926(I19851,g16615);
  not NOT_4927(g19367,I19851);
  not NOT_4928(g19368,g16326);
  not NOT_4929(g19369,g15995);
  not NOT_4930(g19370,g15915);
  not NOT_4931(I19857,g16640);
  not NOT_4932(g19371,I19857);
  not NOT_4933(g19373,g16449);
  not NOT_4934(g19374,g16047);
  not NOT_4935(I19863,g16675);
  not NOT_4936(g19375,I19863);
  not NOT_4937(g19376,g17509);
  not NOT_4938(g19379,g17327);
  not NOT_4939(g19385,g16326);
  not NOT_4940(g19386,g16431);
  not NOT_4941(g19387,g16431);
  not NOT_4942(g19389,g17532);
  not NOT_4943(g19394,g16326);
  not NOT_4944(g19395,g16431);
  not NOT_4945(g19396,g16431);
  not NOT_4946(g19397,g16449);
  not NOT_4947(g19398,g16489);
  not NOT_4948(g19399,g16489);
  not NOT_4949(g19407,g16268);
  not NOT_4950(g19408,g16066);
  not NOT_4951(g19409,g16431);
  not NOT_4952(g19410,g16449);
  not NOT_4953(g19411,g16489);
  not NOT_4954(g19412,g16489);
  not NOT_4955(g19414,g16349);
  not NOT_4956(g19415,g15758);
  not NOT_4957(g19416,g15885);
  not NOT_4958(g19417,g17178);
  not NOT_4959(g19421,g16326);
  not NOT_4960(g19427,g16292);
  not NOT_4961(g19428,g16090);
  not NOT_4962(g19429,g16489);
  not NOT_4963(g19431,g16249);
  not NOT_4964(g19432,g15885);
  not NOT_4965(g19433,g15915);
  not NOT_4966(g19434,g16326);
  not NOT_4967(g19435,g16449);
  not NOT_4968(g19437,g16349);
  not NOT_4969(g19438,g16249);
  not NOT_4970(g19439,g15885);
  not NOT_4971(g19440,g15915);
  not NOT_4972(g19443,g16449);
  not NOT_4973(g19445,g15915);
  not NOT_4974(I19917,g18088);
  not NOT_4975(g19446,I19917);
  not NOT_4976(g19451,g15938);
  not NOT_4977(g19452,g16326);
  not NOT_4978(g19454,g16349);
  not NOT_4979(I19927,g17408);
  not NOT_4980(g19458,I19927);
  not NOT_4981(g19468,g15938);
  not NOT_4982(g19469,g16326);
  not NOT_4983(g19470,g16000);
  not NOT_4984(g19471,g16449);
  not NOT_4985(g19472,g16349);
  not NOT_4986(g19473,g16349);
  not NOT_4987(g19476,g16326);
  not NOT_4988(g19477,g16431);
  not NOT_4989(g19478,g16000);
  not NOT_4990(g19479,g16449);
  not NOT_4991(g19480,g16349);
  not NOT_4992(g19481,g16349);
  not NOT_4993(g19482,g16349);
  not NOT_4994(g19489,g16449);
  not NOT_4995(g19490,g16489);
  not NOT_4996(g19491,g16349);
  not NOT_4997(g19492,g16349);
  not NOT_4998(g19493,g16349);
  not NOT_4999(g19494,g16349);
  not NOT_5000(g19498,g16752);
  not NOT_5001(g19499,g16782);
  not NOT_5002(g19502,g15674);
  not NOT_5003(g19503,g16349);
  not NOT_5004(g19504,g16349);
  not NOT_5005(g19505,g16349);
  not NOT_5006(g19517,g16777);
  not NOT_5007(g19518,g16239);
  not NOT_5008(g19519,g16795);
  not NOT_5009(g19520,g16826);
  not NOT_5010(g19523,g16100);
  not NOT_5011(g19524,g15695);
  not NOT_5012(g19526,g16349);
  not NOT_5013(g19527,g16349);
  not NOT_5014(g19528,g16349);
  not NOT_5015(g19529,g16349);
  not NOT_5016(g19531,g16816);
  not NOT_5017(g19532,g16821);
  not NOT_5018(g19533,g16261);
  not NOT_5019(g19537,g15938);
  not NOT_5020(g19538,g16100);
  not NOT_5021(g19539,g16129);
  not NOT_5022(g19541,g16136);
  not NOT_5023(g19542,g16349);
  not NOT_5024(g19543,g16349);
  not NOT_5025(g19544,g16349);
  not NOT_5026(g19552,g16856);
  not NOT_5027(g19553,g16782);
  not NOT_5028(g19554,g16861);
  not NOT_5029(g19558,g15938);
  not NOT_5030(g19559,g16129);
  not NOT_5031(g19565,g16000);
  not NOT_5032(g19566,g16136);
  not NOT_5033(g19567,g16164);
  not NOT_5034(g19569,g16349);
  not NOT_5035(g19570,g16349);
  not NOT_5036(g19573,g16877);
  not NOT_5037(g19574,g16826);
  not NOT_5038(g19577,g16129);
  not NOT_5039(g19579,g16000);
  not NOT_5040(g19580,g16164);
  not NOT_5041(g19586,g16349);
  not NOT_5042(I20035,g15706);
  not NOT_5043(g19592,I20035);
  not NOT_5044(g19600,g16164);
  not NOT_5045(g19602,g16349);
  not NOT_5046(g19603,g16349);
  not NOT_5047(g19606,g17614);
  not NOT_5048(g19609,g16264);
  not NOT_5049(g19612,g16897);
  not NOT_5050(g19617,g16349);
  not NOT_5051(g19618,g16349);
  not NOT_5052(g19620,g17296);
  not NOT_5053(g19626,g17409);
  not NOT_5054(g19629,g17015);
  not NOT_5055(g19630,g16897);
  not NOT_5056(g19633,g16931);
  not NOT_5057(g19634,g16349);
  not NOT_5058(g19635,g16349);
  not NOT_5059(g19636,g16987);
  not NOT_5060(g19638,g17324);
  not NOT_5061(g19644,g17953);
  not NOT_5062(g19649,g17015);
  not NOT_5063(g19650,g16971);
  not NOT_5064(g19652,g16897);
  not NOT_5065(g19653,g16897);
  not NOT_5066(g19654,g16931);
  not NOT_5067(g19657,g16349);
  not NOT_5068(g19658,g16987);
  not NOT_5069(g19659,g17062);
  not NOT_5070(g19662,g17432);
  not NOT_5071(g19666,g17188);
  not NOT_5072(g19670,g16897);
  not NOT_5073(g19672,g16931);
  not NOT_5074(g19673,g16931);
  not NOT_5075(g19675,g16987);
  not NOT_5076(g19676,g17062);
  not NOT_5077(g19677,g17096);
  not NOT_5078(g19678,g16752);
  not NOT_5079(g19679,g16782);
  not NOT_5080(g19682,g17015);
  not NOT_5081(g19683,g16931);
  not NOT_5082(g19685,g16987);
  not NOT_5083(g19686,g17062);
  not NOT_5084(g19687,g17096);
  not NOT_5085(g19688,g16777);
  not NOT_5086(g19689,g16795);
  not NOT_5087(g19690,g16826);
  not NOT_5088(g19694,g16429);
  not NOT_5089(g19695,g17015);
  not NOT_5090(g19696,g17015);
  not NOT_5091(g19697,g16886);
  not NOT_5092(g19698,g16971);
  not NOT_5093(I20116,g15737);
  not NOT_5094(g19699,I20116);
  not NOT_5095(g19709,g16987);
  not NOT_5096(g19710,g17059);
  not NOT_5097(g19711,g17062);
  not NOT_5098(g19712,g17096);
  not NOT_5099(g19713,g16816);
  not NOT_5100(g19714,g16821);
  not NOT_5101(g19718,g17015);
  not NOT_5102(g19719,g16897);
  not NOT_5103(I20130,g15748);
  not NOT_5104(g19720,I20130);
  not NOT_5105(g19730,g17062);
  not NOT_5106(g19731,g17093);
  not NOT_5107(g19732,g17096);
  not NOT_5108(g19733,g16856);
  not NOT_5109(g19734,g16861);
  not NOT_5110(g19737,g17015);
  not NOT_5111(g19738,g15992);
  not NOT_5112(g19739,g16931);
  not NOT_5113(g19741,g16987);
  not NOT_5114(g19742,g17096);
  not NOT_5115(g19743,g17125);
  not NOT_5116(g19744,g15885);
  not NOT_5117(g19745,g16877);
  not NOT_5118(g19747,g17015);
  not NOT_5119(g19748,g17015);
  not NOT_5120(g19750,g16326);
  not NOT_5121(g19751,g16044);
  not NOT_5122(g19753,g16987);
  not NOT_5123(g19754,g17062);
  not NOT_5124(g19755,g15915);
  not NOT_5125(g19757,g17224);
  not NOT_5126(g19760,g17015);
  not NOT_5127(g19761,g17015);
  not NOT_5128(g19762,g16326);
  not NOT_5129(g19763,g16431);
  not NOT_5130(g19765,g16897);
  not NOT_5131(g19766,g16449);
  not NOT_5132(g19769,g16987);
  not NOT_5133(g19770,g17062);
  not NOT_5134(g19771,g17096);
  not NOT_5135(g19772,g17183);
  not NOT_5136(g19773,g17615);
  not NOT_5137(g19776,g17015);
  not NOT_5138(g19777,g17015);
  not NOT_5139(g19779,g16431);
  not NOT_5140(g19780,g16449);
  not NOT_5141(g19781,g16489);
  not NOT_5142(g19783,g16931);
  not NOT_5143(g19785,g16987);
  not NOT_5144(g19786,g17062);
  not NOT_5145(g19787,g17096);
  not NOT_5146(g19789,g17015);
  not NOT_5147(g19790,g16971);
  not NOT_5148(g19794,g16489);
  not NOT_5149(g19798,g17200);
  not NOT_5150(g19799,g17062);
  not NOT_5151(g19800,g17096);
  not NOT_5152(I20216,g15862);
  not NOT_5153(g19801,I20216);
  not NOT_5154(g19852,g17015);
  not NOT_5155(g19860,g17226);
  not NOT_5156(g19861,g17096);
  not NOT_5157(I20233,g17487);
  not NOT_5158(g19862,I20233);
  not NOT_5159(g19865,g15885);
  not NOT_5160(g19866,g16540);
  not NOT_5161(g19869,g16540);
  not NOT_5162(g19872,g17015);
  not NOT_5163(g19878,g17271);
  not NOT_5164(g19881,g15915);
  not NOT_5165(g19882,g16540);
  not NOT_5166(g19885,g17249);
  not NOT_5167(g19902,g17200);
  not NOT_5168(g19905,g15885);
  not NOT_5169(g19908,g16540);
  not NOT_5170(g19912,g17328);
  not NOT_5171(g19915,g16349);
  not NOT_5172(g19930,g17200);
  not NOT_5173(g19931,g17200);
  not NOT_5174(g19947,g17226);
  not NOT_5175(g19950,g15885);
  not NOT_5176(g19952,g15915);
  not NOT_5177(g19954,g16540);
  not NOT_5178(g19957,g16540);
  not NOT_5179(g19960,g17433);
  not NOT_5180(g19961,g17328);
  not NOT_5181(g19963,g16326);
  not NOT_5182(g19964,g17200);
  not NOT_5183(g19979,g17226);
  not NOT_5184(g19980,g17226);
  not NOT_5185(g19996,g17271);
  not NOT_5186(g19998,g15915);
  not NOT_5187(g20004,g17249);
  not NOT_5188(g20005,g17433);
  not NOT_5189(g20006,g17328);
  not NOT_5190(g20008,g16449);
  not NOT_5191(g20009,g16349);
  not NOT_5192(g20010,g17226);
  not NOT_5193(g20025,g17271);
  not NOT_5194(g20026,g17271);
  not NOT_5195(g20028,g15371);
  not NOT_5196(g20033,g16579);
  not NOT_5197(g20035,g16430);
  not NOT_5198(g20036,g17433);
  not NOT_5199(g20037,g17328);
  not NOT_5200(g20038,g17328);
  not NOT_5201(g20040,g17271);
  not NOT_5202(g20041,g15569);
  not NOT_5203(g20046,g16540);
  not NOT_5204(I20318,g16920);
  not NOT_5205(g20049,I20318);
  not NOT_5206(I20321,g16920);
  not NOT_5207(g20050,I20321);
  not NOT_5208(g20052,g17533);
  not NOT_5209(g20053,g17328);
  not NOT_5210(g20054,g17328);
  not NOT_5211(g20057,g16349);
  not NOT_5212(g20058,g16782);
  not NOT_5213(g20059,g17302);
  not NOT_5214(g20060,g16540);
  not NOT_5215(g20064,g17533);
  not NOT_5216(g20065,g16846);
  not NOT_5217(g20066,g17433);
  not NOT_5218(g20067,g17328);
  not NOT_5219(g20070,g16173);
  not NOT_5220(g20071,g16826);
  not NOT_5221(g20072,g17384);
  not NOT_5222(g20073,g16540);
  not NOT_5223(g20078,g16846);
  not NOT_5224(g20079,g17328);
  not NOT_5225(g20080,g17328);
  not NOT_5226(g20085,g16187);
  not NOT_5227(I20355,g17613);
  not NOT_5228(g20086,I20355);
  not NOT_5229(g20087,g17249);
  not NOT_5230(g20088,g17533);
  not NOT_5231(g20089,g17533);
  not NOT_5232(g20090,g17433);
  not NOT_5233(g20091,g17328);
  not NOT_5234(g20096,g16782);
  not NOT_5235(g20097,g17691);
  not NOT_5236(I20369,g17690);
  not NOT_5237(g20100,I20369);
  not NOT_5238(g20101,g17533);
  not NOT_5239(g20102,g17533);
  not NOT_5240(g20103,g17433);
  not NOT_5241(g20104,g17433);
  not NOT_5242(g20105,g17433);
  not NOT_5243(g20106,g17328);
  not NOT_5244(g20110,g16897);
  not NOT_5245(g20113,g16826);
  not NOT_5246(I20385,g16194);
  not NOT_5247(g20114,I20385);
  not NOT_5248(I20388,g17724);
  not NOT_5249(g20127,I20388);
  not NOT_5250(g20128,g17533);
  not NOT_5251(g20129,g17328);
  not NOT_5252(g20130,g17328);
  not NOT_5253(g20132,g16931);
  not NOT_5254(I20399,g16205);
  not NOT_5255(g20136,I20399);
  not NOT_5256(g20144,g17533);
  not NOT_5257(g20145,g17533);
  not NOT_5258(g20146,g17533);
  not NOT_5259(g20147,g17328);
  not NOT_5260(g20153,g16782);
  not NOT_5261(I20412,g16213);
  not NOT_5262(g20154,I20412);
  not NOT_5263(g20157,g16886);
  not NOT_5264(g20158,g16971);
  not NOT_5265(g20159,g17533);
  not NOT_5266(g20164,g16826);
  not NOT_5267(g20166,g16886);
  not NOT_5268(g20167,g16971);
  not NOT_5269(g20168,g17533);
  not NOT_5270(I20433,g16234);
  not NOT_5271(g20175,I20433);
  not NOT_5272(g20178,g16971);
  not NOT_5273(g20179,g17249);
  not NOT_5274(g20180,g17533);
  not NOT_5275(g20182,g16897);
  not NOT_5276(I20447,g16244);
  not NOT_5277(g20189,I20447);
  not NOT_5278(g20190,g16971);
  not NOT_5279(g20191,g17821);
  not NOT_5280(g20192,g17268);
  not NOT_5281(g20194,g16897);
  not NOT_5282(g20195,g16931);
  not NOT_5283(g20197,g16987);
  not NOT_5284(g20204,g16578);
  not NOT_5285(g20207,g17015);
  not NOT_5286(g20208,g17533);
  not NOT_5287(g20209,g17821);
  not NOT_5288(g20210,g16897);
  not NOT_5289(g20211,g16931);
  not NOT_5290(g20212,g17194);
  not NOT_5291(g20213,g17062);
  not NOT_5292(I20495,g16283);
  not NOT_5293(g20219,I20495);
  not NOT_5294(g20229,g17015);
  not NOT_5295(I20499,g16224);
  not NOT_5296(g20230,I20499);
  not NOT_5297(g20231,g17821);
  not NOT_5298(g20232,g16931);
  not NOT_5299(g20233,g17873);
  not NOT_5300(g20235,g15277);
  not NOT_5301(g20237,g17213);
  not NOT_5302(g20238,g17096);
  not NOT_5303(g20239,g17128);
  not NOT_5304(g20240,g17847);
  not NOT_5305(g20242,g16308);
  not NOT_5306(g20247,g17015);
  not NOT_5307(g20265,g17821);
  not NOT_5308(g20266,g17873);
  not NOT_5309(g20267,g17955);
  not NOT_5310(g20268,g18008);
  not NOT_5311(g20269,g15844);
  not NOT_5312(g20270,g15277);
  not NOT_5313(g20272,g17239);
  not NOT_5314(g20273,g17128);
  not NOT_5315(g20274,g17847);
  not NOT_5316(g20275,g17929);
  not NOT_5317(g20277,g16487);
  not NOT_5318(I20529,g16309);
  not NOT_5319(g20283,I20529);
  not NOT_5320(g20320,g17015);
  not NOT_5321(g20321,g17821);
  not NOT_5322(g20322,g17873);
  not NOT_5323(g20323,g17873);
  not NOT_5324(g20324,g17955);
  not NOT_5325(g20325,g15171);
  not NOT_5326(g20326,g18008);
  not NOT_5327(g20327,g15224);
  not NOT_5328(g20328,g15867);
  not NOT_5329(g20329,g15277);
  not NOT_5330(I20542,g16508);
  not NOT_5331(g20330,I20542);
  not NOT_5332(g20372,g17847);
  not NOT_5333(g20373,g17929);
  not NOT_5334(g20374,g18065);
  not NOT_5335(g20379,g17821);
  not NOT_5336(g20380,g17955);
  not NOT_5337(g20381,g17955);
  not NOT_5338(g20382,g15171);
  not NOT_5339(g20383,g15373);
  not NOT_5340(g20384,g18008);
  not NOT_5341(g20385,g18008);
  not NOT_5342(g20386,g15224);
  not NOT_5343(g20387,g15426);
  not NOT_5344(g20388,g17297);
  not NOT_5345(g20389,g15277);
  not NOT_5346(I20562,g16525);
  not NOT_5347(g20391,I20562);
  not NOT_5348(g20432,g17847);
  not NOT_5349(g20433,g17929);
  not NOT_5350(g20434,g18065);
  not NOT_5351(g20435,g15348);
  not NOT_5352(I20569,g16486);
  not NOT_5353(g20436,I20569);
  not NOT_5354(g20441,g17873);
  not NOT_5355(g20442,g15171);
  not NOT_5356(g20443,g15171);
  not NOT_5357(g20444,g15373);
  not NOT_5358(g20445,g15224);
  not NOT_5359(g20446,g15224);
  not NOT_5360(g20447,g15426);
  not NOT_5361(g20448,g15509);
  not NOT_5362(g20449,g15277);
  not NOT_5363(g20450,g15277);
  not NOT_5364(g20451,g15277);
  not NOT_5365(g20452,g17200);
  not NOT_5366(I20584,g16587);
  not NOT_5367(g20453,I20584);
  not NOT_5368(g20494,g17847);
  not NOT_5369(g20495,g17926);
  not NOT_5370(g20496,g17929);
  not NOT_5371(g20497,g18065);
  not NOT_5372(g20498,g15348);
  not NOT_5373(g20499,g15483);
  not NOT_5374(g20500,g17873);
  not NOT_5375(g20501,g17955);
  not NOT_5376(g20502,g15373);
  not NOT_5377(g20503,g15373);
  not NOT_5378(g20504,g18008);
  not NOT_5379(g20505,g15426);
  not NOT_5380(g20506,g15426);
  not NOT_5381(g20507,g15509);
  not NOT_5382(g20508,g15277);
  not NOT_5383(g20509,g15277);
  not NOT_5384(g20510,g17226);
  not NOT_5385(g20511,g17929);
  not NOT_5386(g20512,g18062);
  not NOT_5387(g20513,g18065);
  not NOT_5388(g20514,g15348);
  not NOT_5389(g20515,g15483);
  not NOT_5390(I20609,g16539);
  not NOT_5391(g20516,I20609);
  not NOT_5392(g20523,g17821);
  not NOT_5393(g20524,g17873);
  not NOT_5394(g20525,g17955);
  not NOT_5395(g20526,g15171);
  not NOT_5396(g20527,g18008);
  not NOT_5397(g20528,g15224);
  not NOT_5398(g20529,g15509);
  not NOT_5399(g20530,g15509);
  not NOT_5400(g20531,g15907);
  not NOT_5401(g20532,g15277);
  not NOT_5402(g20533,g17271);
  not NOT_5403(g20534,g17183);
  not NOT_5404(g20535,g17847);
  not NOT_5405(g20536,g18065);
  not NOT_5406(g20537,g15345);
  not NOT_5407(g20538,g15348);
  not NOT_5408(g20539,g15483);
  not NOT_5409(g20540,g16646);
  not NOT_5410(g20541,g17821);
  not NOT_5411(g20542,g17873);
  not NOT_5412(g20543,g17955);
  not NOT_5413(g20544,g15171);
  not NOT_5414(g20545,g15373);
  not NOT_5415(g20546,g18008);
  not NOT_5416(g20547,g15224);
  not NOT_5417(g20548,g15426);
  not NOT_5418(g20549,g15277);
  not NOT_5419(g20550,g15864);
  not NOT_5420(g20551,g17302);
  not NOT_5421(g20552,g17847);
  not NOT_5422(g20553,g17929);
  not NOT_5423(g20554,g15348);
  not NOT_5424(g20555,g15480);
  not NOT_5425(g20556,g15483);
  not NOT_5426(I20647,g17010);
  not NOT_5427(g20557,I20647);
  not NOT_5428(I20650,g17010);
  not NOT_5429(g20558,I20650);
  not NOT_5430(g20560,g17328);
  not NOT_5431(g20561,g17873);
  not NOT_5432(g20562,g17955);
  not NOT_5433(g20563,g15171);
  not NOT_5434(g20564,g15373);
  not NOT_5435(g20565,g18008);
  not NOT_5436(g20566,g15224);
  not NOT_5437(g20567,g15426);
  not NOT_5438(g20568,g15509);
  not NOT_5439(g20569,g15277);
  not NOT_5440(g20570,g15277);
  not NOT_5441(g20571,g15277);
  not NOT_5442(g20572,g15833);
  not NOT_5443(g20573,g17384);
  not NOT_5444(g20574,g17847);
  not NOT_5445(g20575,g17929);
  not NOT_5446(g20576,g18065);
  not NOT_5447(g20577,g15483);
  not NOT_5448(g20578,g15563);
  not NOT_5449(g20579,g17249);
  not NOT_5450(g20580,g17328);
  not NOT_5451(g20582,g17873);
  not NOT_5452(g20583,g17873);
  not NOT_5453(g20584,g17873);
  not NOT_5454(g20585,g17955);
  not NOT_5455(g20586,g15171);
  not NOT_5456(g20587,g15373);
  not NOT_5457(g20588,g18008);
  not NOT_5458(g20589,g15224);
  not NOT_5459(g20590,g15426);
  not NOT_5460(g20591,g15509);
  not NOT_5461(g20592,g15277);
  not NOT_5462(g20593,g15277);
  not NOT_5463(g20594,g15277);
  not NOT_5464(g20595,g15877);
  not NOT_5465(I20690,g15733);
  not NOT_5466(g20596,I20690);
  not NOT_5467(g20597,g17847);
  not NOT_5468(g20598,g17929);
  not NOT_5469(g20599,g18065);
  not NOT_5470(g20600,g15348);
  not NOT_5471(g20601,g17433);
  not NOT_5472(g20603,g17873);
  not NOT_5473(g20604,g17873);
  not NOT_5474(g20605,g17955);
  not NOT_5475(g20606,g17955);
  not NOT_5476(g20607,g17955);
  not NOT_5477(g20608,g15171);
  not NOT_5478(g20609,g15373);
  not NOT_5479(g20610,g18008);
  not NOT_5480(g20611,g18008);
  not NOT_5481(g20612,g18008);
  not NOT_5482(g20613,g15224);
  not NOT_5483(g20614,g15426);
  not NOT_5484(g20615,g15509);
  not NOT_5485(g20616,g15277);
  not NOT_5486(g20617,g15277);
  not NOT_5487(g20618,g15277);
  not NOT_5488(g20622,g15595);
  not NOT_5489(g20623,g17929);
  not NOT_5490(g20624,g18065);
  not NOT_5491(g20625,g15348);
  not NOT_5492(g20626,g15483);
  not NOT_5493(g20627,g17433);
  not NOT_5494(g20629,g17955);
  not NOT_5495(g20630,g17955);
  not NOT_5496(g20631,g15171);
  not NOT_5497(g20632,g15171);
  not NOT_5498(g20633,g15171);
  not NOT_5499(g20634,g15373);
  not NOT_5500(g20635,g18008);
  not NOT_5501(g20636,g18008);
  not NOT_5502(g20637,g15224);
  not NOT_5503(g20638,g15224);
  not NOT_5504(g20639,g15224);
  not NOT_5505(g20640,g15426);
  not NOT_5506(g20641,g15509);
  not NOT_5507(g20642,g15277);
  not NOT_5508(g20643,g15962);
  not NOT_5509(g20648,g15615);
  not NOT_5510(g20649,g18065);
  not NOT_5511(g20650,g15348);
  not NOT_5512(g20651,g15483);
  not NOT_5513(I20744,g17141);
  not NOT_5514(g20652,I20744);
  not NOT_5515(I20747,g17141);
  not NOT_5516(g20653,I20747);
  not NOT_5517(I20750,g16677);
  not NOT_5518(g20654,I20750);
  not NOT_5519(I20753,g16677);
  not NOT_5520(g20655,I20753);
  not NOT_5521(g20656,g17249);
  not NOT_5522(g20657,g17433);
  not NOT_5523(g20659,g17873);
  not NOT_5524(g20660,g17873);
  not NOT_5525(g20661,g15171);
  not NOT_5526(g20662,g15171);
  not NOT_5527(g20663,g15373);
  not NOT_5528(g20664,g15373);
  not NOT_5529(g20665,g15373);
  not NOT_5530(g20666,g15224);
  not NOT_5531(g20667,g15224);
  not NOT_5532(g20668,g15426);
  not NOT_5533(g20669,g15426);
  not NOT_5534(g20670,g15426);
  not NOT_5535(g20671,g15509);
  not NOT_5536(g20672,g15277);
  not NOT_5537(g20673,g15277);
  not NOT_5538(g20674,g15277);
  not NOT_5539(g20679,g15634);
  not NOT_5540(g20680,g15348);
  not NOT_5541(g20681,g15483);
  not NOT_5542(I20781,g17155);
  not NOT_5543(g20695,I20781);
  not NOT_5544(g20696,g17533);
  not NOT_5545(g20697,g17433);
  not NOT_5546(g20698,g17873);
  not NOT_5547(g20699,g17873);
  not NOT_5548(g20700,g17873);
  not NOT_5549(g20701,g17955);
  not NOT_5550(g20702,g17955);
  not NOT_5551(g20703,g15373);
  not NOT_5552(g20704,g15373);
  not NOT_5553(I20793,g17694);
  not NOT_5554(g20705,I20793);
  not NOT_5555(g20706,g18008);
  not NOT_5556(g20707,g18008);
  not NOT_5557(g20708,g15426);
  not NOT_5558(g20709,g15426);
  not NOT_5559(g20710,g15509);
  not NOT_5560(g20711,g15509);
  not NOT_5561(g20712,g15509);
  not NOT_5562(g20713,g15277);
  not NOT_5563(g20714,g15277);
  not NOT_5564(g20715,g15277);
  not NOT_5565(g20716,g15277);
  not NOT_5566(g20732,g15595);
  not NOT_5567(g20737,g15656);
  not NOT_5568(g20738,g15483);
  not NOT_5569(I20816,g17088);
  not NOT_5570(g20763,I20816);
  not NOT_5571(I20819,g17088);
  not NOT_5572(g20764,I20819);
  not NOT_5573(g20765,g17748);
  not NOT_5574(g20766,g17433);
  not NOT_5575(g20767,g17873);
  not NOT_5576(g20768,g17955);
  not NOT_5577(g20769,g17955);
  not NOT_5578(g20770,g17955);
  not NOT_5579(g20771,g15171);
  not NOT_5580(g20772,g15171);
  not NOT_5581(I20830,g17657);
  not NOT_5582(g20773,I20830);
  not NOT_5583(g20774,g18008);
  not NOT_5584(g20775,g18008);
  not NOT_5585(g20776,g18008);
  not NOT_5586(g20777,g15224);
  not NOT_5587(g20778,g15224);
  not NOT_5588(g20779,g15509);
  not NOT_5589(g20780,g15509);
  not NOT_5590(I20840,g17727);
  not NOT_5591(g20781,I20840);
  not NOT_5592(g20782,g15853);
  not NOT_5593(I20846,g16923);
  not NOT_5594(g20785,I20846);
  not NOT_5595(g20852,g15595);
  not NOT_5596(g20853,g15595);
  not NOT_5597(g20869,g15615);
  not NOT_5598(g20874,g15680);
  not NOT_5599(I20861,g16960);
  not NOT_5600(g20899,I20861);
  not NOT_5601(I20864,g16960);
  not NOT_5602(g20900,I20864);
  not NOT_5603(I20867,g16216);
  not NOT_5604(g20901,I20867);
  not NOT_5605(I20870,g16216);
  not NOT_5606(g20902,I20870);
  not NOT_5607(g20903,g17249);
  not NOT_5608(g20904,g17433);
  not NOT_5609(g20909,g17955);
  not NOT_5610(g20910,g15171);
  not NOT_5611(g20911,g15171);
  not NOT_5612(g20912,g15171);
  not NOT_5613(g20913,g15373);
  not NOT_5614(g20914,g15373);
  not NOT_5615(I20882,g17619);
  not NOT_5616(g20915,I20882);
  not NOT_5617(g20916,g18008);
  not NOT_5618(g20917,g15224);
  not NOT_5619(g20918,g15224);
  not NOT_5620(g20919,g15224);
  not NOT_5621(g20920,g15426);
  not NOT_5622(g20921,g15426);
  not NOT_5623(I20891,g17700);
  not NOT_5624(g20922,I20891);
  not NOT_5625(g20923,g15277);
  not NOT_5626(I20895,g16954);
  not NOT_5627(g20924,I20895);
  not NOT_5628(g20978,g15595);
  not NOT_5629(g20993,g15615);
  not NOT_5630(g20994,g15615);
  not NOT_5631(g21010,g15634);
  not NOT_5632(I20910,g17197);
  not NOT_5633(g21036,I20910);
  not NOT_5634(I20913,g16964);
  not NOT_5635(g21037,I20913);
  not NOT_5636(g21048,g17533);
  not NOT_5637(g21049,g17433);
  not NOT_5638(g21050,g17873);
  not NOT_5639(g21051,g15171);
  not NOT_5640(g21052,g15373);
  not NOT_5641(g21053,g15373);
  not NOT_5642(g21054,g15373);
  not NOT_5643(g21055,g15224);
  not NOT_5644(g21056,g15426);
  not NOT_5645(g21057,g15426);
  not NOT_5646(g21058,g15426);
  not NOT_5647(g21059,g15509);
  not NOT_5648(g21060,g15509);
  not NOT_5649(I20929,g17663);
  not NOT_5650(g21061,I20929);
  not NOT_5651(g21068,g15277);
  not NOT_5652(g21069,g15277);
  not NOT_5653(I20937,g16967);
  not NOT_5654(g21070,I20937);
  not NOT_5655(g21123,g15615);
  not NOT_5656(g21138,g15634);
  not NOT_5657(g21139,g15634);
  not NOT_5658(g21155,g15656);
  not NOT_5659(g21156,g17247);
  not NOT_5660(g21160,g17508);
  not NOT_5661(I20951,g17782);
  not NOT_5662(g21175,I20951);
  not NOT_5663(I20954,g16228);
  not NOT_5664(g21176,I20954);
  not NOT_5665(I20957,g16228);
  not NOT_5666(g21177,I20957);
  not NOT_5667(g21178,g17955);
  not NOT_5668(g21179,g15373);
  not NOT_5669(g21180,g18008);
  not NOT_5670(g21181,g15426);
  not NOT_5671(g21182,g15509);
  not NOT_5672(g21183,g15509);
  not NOT_5673(g21184,g15509);
  not NOT_5674(g21185,g15277);
  not NOT_5675(g21189,g15634);
  not NOT_5676(g21204,g15656);
  not NOT_5677(g21205,g15656);
  not NOT_5678(g21221,g15680);
  not NOT_5679(g21222,g17430);
  not NOT_5680(g21225,g17428);
  not NOT_5681(g21228,g17531);
  not NOT_5682(I20982,g16300);
  not NOT_5683(g21245,I20982);
  not NOT_5684(I20985,g16300);
  not NOT_5685(g21246,I20985);
  not NOT_5686(g21247,g15171);
  not NOT_5687(g21248,g15224);
  not NOT_5688(g21249,g15509);
  not NOT_5689(g21252,g15656);
  not NOT_5690(g21267,g15680);
  not NOT_5691(g21268,g15680);
  not NOT_5692(g21269,g15506);
  not NOT_5693(I20999,g16709);
  not NOT_5694(g21270,I20999);
  not NOT_5695(I21002,g16709);
  not NOT_5696(g21271,I21002);
  not NOT_5697(I21006,g15579);
  not NOT_5698(g21273,I21006);
  not NOT_5699(g21274,g15373);
  not NOT_5700(g21275,g15426);
  not NOT_5701(I21013,g15806);
  not NOT_5702(g21278,I21013);
  not NOT_5703(g21279,g15680);
  not NOT_5704(g21280,g16601);
  not NOT_5705(g21281,g16286);
  not NOT_5706(I21019,g17325);
  not NOT_5707(g21282,I21019);
  not NOT_5708(g21286,g15509);
  not NOT_5709(I21029,g15816);
  not NOT_5710(g21290,I21029);
  not NOT_5711(g21291,g16620);
  not NOT_5712(I21033,g17221);
  not NOT_5713(g21292,I21033);
  not NOT_5714(I21036,g17221);
  not NOT_5715(g21293,I21036);
  not NOT_5716(g21295,g17533);
  not NOT_5717(I21042,g15824);
  not NOT_5718(g21297,I21042);
  not NOT_5719(g21299,g16600);
  not NOT_5720(I21047,g17429);
  not NOT_5721(g21300,I21047);
  not NOT_5722(g21304,g17367);
  not NOT_5723(g21305,g15758);
  not NOT_5724(g21306,g15582);
  not NOT_5725(g21308,g17485);
  not NOT_5726(I21058,g17747);
  not NOT_5727(g21326,I21058);
  not NOT_5728(g21329,g16577);
  not NOT_5729(I21067,g15573);
  not NOT_5730(g21335,I21067);
  not NOT_5731(g21336,g17367);
  not NOT_5732(g21337,g15758);
  not NOT_5733(I21074,g17766);
  not NOT_5734(g21340,I21074);
  not NOT_5735(g21343,g16428);
  not NOT_5736(g21346,g17821);
  not NOT_5737(g21349,g15758);
  not NOT_5738(g21352,g16322);
  not NOT_5739(g21355,g17821);
  not NOT_5740(g21358,g16307);
  not NOT_5741(g21362,g17873);
  not NOT_5742(I21100,g16284);
  not NOT_5743(g21366,I21100);
  not NOT_5744(g21369,g16285);
  not NOT_5745(g21370,g16323);
  not NOT_5746(g21379,g17873);
  not NOT_5747(g21380,g17955);
  not NOT_5748(g21381,g18008);
  not NOT_5749(g21383,g17367);
  not NOT_5750(I21115,g15714);
  not NOT_5751(g21387,I21115);
  not NOT_5752(g21393,g17264);
  not NOT_5753(g21395,g17873);
  not NOT_5754(g21396,g17955);
  not NOT_5755(g21397,g15171);
  not NOT_5756(g21398,g18008);
  not NOT_5757(g21399,g15224);
  not NOT_5758(g21400,g17847);
  not NOT_5759(g21406,g17955);
  not NOT_5760(g21407,g15171);
  not NOT_5761(g21408,g15373);
  not NOT_5762(g21409,g18008);
  not NOT_5763(g21410,g15224);
  not NOT_5764(g21411,g15426);
  not NOT_5765(g21412,g15758);
  not NOT_5766(g21413,g15585);
  not NOT_5767(g21414,g17929);
  not NOT_5768(g21418,g17821);
  not NOT_5769(g21421,g15171);
  not NOT_5770(g21422,g15373);
  not NOT_5771(g21423,g15224);
  not NOT_5772(g21424,g15426);
  not NOT_5773(g21425,g15509);
  not NOT_5774(g21426,g15277);
  not NOT_5775(g21427,g17367);
  not NOT_5776(g21428,g15758);
  not NOT_5777(g21430,g15608);
  not NOT_5778(g21431,g18065);
  not NOT_5779(g21434,g17248);
  not NOT_5780(I21162,g17292);
  not NOT_5781(g21451,I21162);
  not NOT_5782(g21454,g15373);
  not NOT_5783(g21455,g15426);
  not NOT_5784(g21456,g15509);
  not NOT_5785(g21457,g17367);
  not NOT_5786(g21458,g15758);
  not NOT_5787(g21460,g15628);
  not NOT_5788(g21461,g15348);
  not NOT_5789(g21463,g15588);
  not NOT_5790(g21466,g15509);
  not NOT_5791(g21467,g15758);
  not NOT_5792(I21181,g17413);
  not NOT_5793(g21468,I21181);
  not NOT_5794(g21510,g15647);
  not NOT_5795(g21511,g15483);
  not NOT_5796(I21189,g17475);
  not NOT_5797(g21514,I21189);
  not NOT_5798(g21556,g15669);
  not NOT_5799(g21560,g17873);
  not NOT_5800(g21561,g15595);
  not NOT_5801(I21199,g17501);
  not NOT_5802(g21562,I21199);
  not NOT_5803(g21604,g15938);
  not NOT_5804(g21607,g17873);
  not NOT_5805(g21608,g17955);
  not NOT_5806(g21609,g18008);
  not NOT_5807(g21610,g15615);
  not NOT_5808(I21210,g17526);
  not NOT_5809(g21611,I21210);
  not NOT_5810(g21653,g17663);
  not NOT_5811(g21654,g17619);
  not NOT_5812(g21656,g17700);
  not NOT_5813(g21657,g17657);
  not NOT_5814(g21659,g17727);
  not NOT_5815(g21660,g17694);
  not NOT_5816(I21222,g18091);
  not NOT_5817(g21661,I21222);
  not NOT_5818(g21662,g16540);
  not NOT_5819(I21226,g16540);
  not NOT_5820(g21665,I21226);
  not NOT_5821(g21666,g16540);
  not NOT_5822(I21230,g16540);
  not NOT_5823(g21669,I21230);
  not NOT_5824(g21670,g16540);
  not NOT_5825(I21234,g16540);
  not NOT_5826(g21673,I21234);
  not NOT_5827(g21674,g16540);
  not NOT_5828(I21238,g16540);
  not NOT_5829(g21677,I21238);
  not NOT_5830(g21678,g16540);
  not NOT_5831(I21242,g16540);
  not NOT_5832(g21681,I21242);
  not NOT_5833(g21682,g16540);
  not NOT_5834(I21246,g16540);
  not NOT_5835(g21685,I21246);
  not NOT_5836(g21686,g16540);
  not NOT_5837(I21250,g16540);
  not NOT_5838(g21689,I21250);
  not NOT_5839(g21690,g16540);
  not NOT_5840(I21254,g16540);
  not NOT_5841(g21693,I21254);
  not NOT_5842(g21694,g16540);
  not NOT_5843(I21258,g16540);
  not NOT_5844(g21697,I21258);
  not NOT_5845(g21698,g18562);
  not NOT_5846(I21285,g18215);
  not NOT_5847(g21722,I21285);
  not NOT_5848(I21288,g18216);
  not NOT_5849(g21723,I21288);
  not NOT_5850(I21291,g18273);
  not NOT_5851(g21724,I21291);
  not NOT_5852(I21294,g18274);
  not NOT_5853(g21725,I21294);
  not NOT_5854(I21297,g18597);
  not NOT_5855(g21726,I21297);
  not NOT_5856(I21300,g18598);
  not NOT_5857(g21727,I21300);
  not NOT_5858(I21477,g18695);
  not NOT_5859(g21902,I21477);
  not NOT_5860(I21480,g18696);
  not NOT_5861(g21903,I21480);
  not NOT_5862(I21483,g18726);
  not NOT_5863(g21904,I21483);
  not NOT_5864(I21486,g18727);
  not NOT_5865(g21905,I21486);
  not NOT_5866(g22136,g20277);
  not NOT_5867(g22137,g21370);
  not NOT_5868(g22138,g21370);
  not NOT_5869(I21722,g19264);
  not NOT_5870(g22139,I21722);
  not NOT_5871(g22144,g18997);
  not NOT_5872(g22146,g18997);
  not NOT_5873(g22147,g18997);
  not NOT_5874(g22148,g19074);
  not NOT_5875(g22150,g21280);
  not NOT_5876(I21734,g19268);
  not NOT_5877(g22151,I21734);
  not NOT_5878(g22153,g18997);
  not NOT_5879(g22154,g19074);
  not NOT_5880(g22155,g19074);
  not NOT_5881(g22156,g19147);
  not NOT_5882(I21744,g19338);
  not NOT_5883(g22159,I21744);
  not NOT_5884(g22166,g18997);
  not NOT_5885(g22167,g19074);
  not NOT_5886(g22168,g19147);
  not NOT_5887(g22169,g19147);
  not NOT_5888(g22170,g19210);
  not NOT_5889(g22171,g18882);
  not NOT_5890(I21757,g21308);
  not NOT_5891(g22173,I21757);
  not NOT_5892(g22176,g18997);
  not NOT_5893(g22177,g19074);
  not NOT_5894(g22178,g19147);
  not NOT_5895(g22179,g19210);
  not NOT_5896(g22180,g19210);
  not NOT_5897(g22181,g19277);
  not NOT_5898(I21766,g19620);
  not NOT_5899(g22182,I21766);
  not NOT_5900(I21769,g19402);
  not NOT_5901(g22189,I21769);
  not NOT_5902(g22192,g19801);
  not NOT_5903(I21776,g21308);
  not NOT_5904(g22194,I21776);
  not NOT_5905(g22197,g19074);
  not NOT_5906(g22198,g19147);
  not NOT_5907(g22199,g19210);
  not NOT_5908(g22200,g19277);
  not NOT_5909(g22201,g19277);
  not NOT_5910(I21784,g19638);
  not NOT_5911(g22202,I21784);
  not NOT_5912(I21787,g19422);
  not NOT_5913(g22207,I21787);
  not NOT_5914(I21792,g21308);
  not NOT_5915(g22210,I21792);
  not NOT_5916(g22213,g19147);
  not NOT_5917(g22214,g19210);
  not NOT_5918(g22215,g19277);
  not NOT_5919(I21802,g21308);
  not NOT_5920(g22220,I21802);
  not NOT_5921(g22223,g19210);
  not NOT_5922(g22224,g19277);
  not NOT_5923(g22227,g19801);
  not NOT_5924(I21810,g20596);
  not NOT_5925(g22228,I21810);
  not NOT_5926(I21815,g21308);
  not NOT_5927(g22300,I21815);
  not NOT_5928(g22303,g19277);
  not NOT_5929(g22305,g19801);
  not NOT_5930(g22311,g18935);
  not NOT_5931(g22317,g19801);
  not NOT_5932(I21831,g19127);
  not NOT_5933(g22319,I21831);
  not NOT_5934(g22330,g19801);
  not NOT_5935(I21838,g19263);
  not NOT_5936(g22332,I21838);
  not NOT_5937(g22338,g19801);
  not NOT_5938(g22339,g19801);
  not NOT_5939(g22341,g19801);
  not NOT_5940(g22358,g19801);
  not NOT_5941(g22359,g19495);
  not NOT_5942(I21849,g19620);
  not NOT_5943(g22360,I21849);
  not NOT_5944(g22406,g19506);
  not NOT_5945(g22407,g19455);
  not NOT_5946(g22408,g19483);
  not NOT_5947(I21860,g19638);
  not NOT_5948(g22409,I21860);
  not NOT_5949(g22449,g19597);
  not NOT_5950(g22455,g19801);
  not NOT_5951(g22456,g19801);
  not NOT_5952(g22492,g19614);
  not NOT_5953(g22493,g19801);
  not NOT_5954(g22494,g19801);
  not NOT_5955(g22495,g19801);
  not NOT_5956(g22496,g19510);
  not NOT_5957(g22497,g19513);
  not NOT_5958(g22519,g19801);
  not NOT_5959(g22520,g19801);
  not NOT_5960(g22526,g19801);
  not NOT_5961(g22527,g19546);
  not NOT_5962(g22528,g19801);
  not NOT_5963(g22529,g19549);
  not NOT_5964(I21911,g21278);
  not NOT_5965(g22541,I21911);
  not NOT_5966(g22542,g19801);
  not NOT_5967(g22543,g19801);
  not NOT_5968(g22544,g19589);
  not NOT_5969(I21918,g21290);
  not NOT_5970(g22546,I21918);
  not NOT_5971(I21922,g21335);
  not NOT_5972(g22550,I21922);
  not NOT_5973(I21930,g21297);
  not NOT_5974(g22592,I21930);
  not NOT_5975(g22593,g19801);
  not NOT_5976(I21934,g21273);
  not NOT_5977(g22594,I21934);
  not NOT_5978(I21941,g18918);
  not NOT_5979(g22626,I21941);
  not NOT_5980(g22635,g19801);
  not NOT_5981(g22646,g19389);
  not NOT_5982(I21959,g20242);
  not NOT_5983(g22647,I21959);
  not NOT_5984(g22649,g19063);
  not NOT_5985(I21969,g21370);
  not NOT_5986(g22658,I21969);
  not NOT_5987(g22660,g19140);
  not NOT_5988(g22667,g21156);
  not NOT_5989(g22682,g19379);
  not NOT_5990(I22000,g20277);
  not NOT_5991(g22683,I22000);
  not NOT_5992(I22009,g21269);
  not NOT_5993(g22698,I22009);
  not NOT_5994(g22714,g20436);
  not NOT_5995(g22716,g19795);
  not NOT_5996(g22718,g20887);
  not NOT_5997(I22024,g19350);
  not NOT_5998(g22719,I22024);
  not NOT_5999(I22028,g20204);
  not NOT_6000(g22721,I22028);
  not NOT_6001(I22031,g21387);
  not NOT_6002(g22722,I22031);
  not NOT_6003(g22756,g20436);
  not NOT_6004(g22758,g20330);
  not NOT_6005(g22759,g19857);
  not NOT_6006(g22761,g21024);
  not NOT_6007(I22046,g19330);
  not NOT_6008(g22763,I22046);
  not NOT_6009(g22830,g20283);
  not NOT_6010(g22840,g20330);
  not NOT_6011(g22841,g20391);
  not NOT_6012(g22842,g19875);
  not NOT_6013(g22844,g21163);
  not NOT_6014(g22845,g20682);
  not NOT_6015(g22847,g20283);
  not NOT_6016(g22854,g20330);
  not NOT_6017(g22855,g20391);
  not NOT_6018(g22856,g20453);
  not NOT_6019(g22857,g20739);
  not NOT_6020(g22858,g20751);
  not NOT_6021(g22860,g20000);
  not NOT_6022(g22865,g20330);
  not NOT_6023(g22866,g20330);
  not NOT_6024(g22867,g20391);
  not NOT_6025(g22868,g20453);
  not NOT_6026(g22869,g20875);
  not NOT_6027(g22870,g20887);
  not NOT_6028(I22096,g19890);
  not NOT_6029(g22881,I22096);
  not NOT_6030(g22882,g20391);
  not NOT_6031(g22883,g20391);
  not NOT_6032(g22884,g20453);
  not NOT_6033(g22896,g21012);
  not NOT_6034(g22897,g21024);
  not NOT_6035(g22898,g20283);
  not NOT_6036(g22903,g20330);
  not NOT_6037(I22111,g19919);
  not NOT_6038(g22904,I22111);
  not NOT_6039(I22114,g19935);
  not NOT_6040(g22905,I22114);
  not NOT_6041(g22906,g20453);
  not NOT_6042(g22907,g20453);
  not NOT_6043(g22919,g21163);
  not NOT_6044(g22922,g20330);
  not NOT_6045(I22124,g21300);
  not NOT_6046(g22923,I22124);
  not NOT_6047(g22926,g20391);
  not NOT_6048(I22128,g19968);
  not NOT_6049(g22927,I22128);
  not NOT_6050(I22131,g19984);
  not NOT_6051(g22928,I22131);
  not NOT_6052(g22935,g20283);
  not NOT_6053(g22936,g20283);
  not NOT_6054(I22143,g20189);
  not NOT_6055(g22957,I22143);
  not NOT_6056(g22973,g20330);
  not NOT_6057(g22974,g20330);
  not NOT_6058(g22975,g20391);
  not NOT_6059(I22149,g21036);
  not NOT_6060(g22976,I22149);
  not NOT_6061(g22979,g20453);
  not NOT_6062(I22153,g20014);
  not NOT_6063(g22980,I22153);
  not NOT_6064(g22981,g20283);
  not NOT_6065(g22985,g20330);
  not NOT_6066(g22986,g20330);
  not NOT_6067(g22987,g20391);
  not NOT_6068(g22988,g20391);
  not NOT_6069(g22989,g20453);
  not NOT_6070(g22994,g20436);
  not NOT_6071(g22995,g20330);
  not NOT_6072(g22996,g20330);
  not NOT_6073(g22997,g20391);
  not NOT_6074(g22998,g20391);
  not NOT_6075(g22999,g20453);
  not NOT_6076(g23000,g20453);
  not NOT_6077(g23001,g19801);
  not NOT_6078(I22177,g21366);
  not NOT_6079(g23002,I22177);
  not NOT_6080(I22180,g21366);
  not NOT_6081(g23003,I22180);
  not NOT_6082(g23004,g20283);
  not NOT_6083(g23005,g20283);
  not NOT_6084(g23011,g20330);
  not NOT_6085(g23012,g20330);
  not NOT_6086(g23013,g20330);
  not NOT_6087(g23014,g20391);
  not NOT_6088(g23015,g20391);
  not NOT_6089(g23016,g20453);
  not NOT_6090(g23017,g20453);
  not NOT_6091(g23018,g19801);
  not NOT_6092(g23019,g19866);
  not NOT_6093(g23020,g19869);
  not NOT_6094(g23021,g20283);
  not NOT_6095(g23022,g20283);
  not NOT_6096(g23026,g20391);
  not NOT_6097(g23027,g20391);
  not NOT_6098(g23028,g20391);
  not NOT_6099(g23029,g20453);
  not NOT_6100(g23030,g20453);
  not NOT_6101(g23031,g19801);
  not NOT_6102(I22211,g21463);
  not NOT_6103(g23032,I22211);
  not NOT_6104(g23041,g19882);
  not NOT_6105(g23046,g20283);
  not NOT_6106(g23055,g20887);
  not NOT_6107(g23057,g20453);
  not NOT_6108(g23058,g20453);
  not NOT_6109(g23059,g20453);
  not NOT_6110(g23060,g19908);
  not NOT_6111(g23061,g20283);
  not NOT_6112(g23066,g20330);
  not NOT_6113(g23082,g21024);
  not NOT_6114(g23084,g19954);
  not NOT_6115(g23085,g19957);
  not NOT_6116(g23086,g20283);
  not NOT_6117(I22240,g20086);
  not NOT_6118(g23088,I22240);
  not NOT_6119(g23111,g20391);
  not NOT_6120(g23127,g21163);
  not NOT_6121(g23128,g20283);
  not NOT_6122(g23138,g20453);
  not NOT_6123(g23152,g20283);
  not NOT_6124(I22264,g20100);
  not NOT_6125(g23154,I22264);
  not NOT_6126(g23170,g20046);
  not NOT_6127(I22275,g20127);
  not NOT_6128(g23172,I22275);
  not NOT_6129(g23182,g21389);
  not NOT_6130(g23189,g20060);
  not NOT_6131(I22286,g19446);
  not NOT_6132(g23190,I22286);
  not NOT_6133(I22289,g19446);
  not NOT_6134(g23191,I22289);
  not NOT_6135(g23192,g20248);
  not NOT_6136(g23196,g20785);
  not NOT_6137(I22302,g19353);
  not NOT_6138(g23202,I22302);
  not NOT_6139(g23203,g20073);
  not NOT_6140(g23211,g21308);
  not NOT_6141(g23214,g20785);
  not NOT_6142(g23215,g20785);
  not NOT_6143(g23216,g20924);
  not NOT_6144(I22316,g19361);
  not NOT_6145(g23219,I22316);
  not NOT_6146(g23221,g20785);
  not NOT_6147(g23222,g20785);
  not NOT_6148(g23223,g21308);
  not NOT_6149(g23226,g20924);
  not NOT_6150(g23227,g20924);
  not NOT_6151(g23228,g21070);
  not NOT_6152(I22327,g19367);
  not NOT_6153(g23230,I22327);
  not NOT_6154(g23231,g20050);
  not NOT_6155(I22331,g19417);
  not NOT_6156(g23232,I22331);
  not NOT_6157(g23233,g21037);
  not NOT_6158(g23234,g20375);
  not NOT_6159(g23235,g20785);
  not NOT_6160(g23236,g20785);
  not NOT_6161(g23237,g20924);
  not NOT_6162(g23238,g20924);
  not NOT_6163(g23239,g21308);
  not NOT_6164(g23242,g21070);
  not NOT_6165(g23243,g21070);
  not NOT_6166(I22343,g19371);
  not NOT_6167(g23244,I22343);
  not NOT_6168(g23245,g20785);
  not NOT_6169(g23246,g20785);
  not NOT_6170(g23247,g20924);
  not NOT_6171(g23248,g20924);
  not NOT_6172(g23249,g21070);
  not NOT_6173(g23250,g21070);
  not NOT_6174(I22353,g19375);
  not NOT_6175(g23252,I22353);
  not NOT_6176(g23253,g21037);
  not NOT_6177(g23256,g20785);
  not NOT_6178(g23257,g20924);
  not NOT_6179(g23258,g20924);
  not NOT_6180(g23259,g21070);
  not NOT_6181(g23260,g21070);
  not NOT_6182(I22366,g19757);
  not NOT_6183(g23263,I22366);
  not NOT_6184(g23264,g21037);
  not NOT_6185(g23267,g20097);
  not NOT_6186(g23270,g20785);
  not NOT_6187(g23271,g20785);
  not NOT_6188(g23272,g20924);
  not NOT_6189(g23273,g21070);
  not NOT_6190(g23274,g21070);
  not NOT_6191(I22380,g21156);
  not NOT_6192(g23277,I22380);
  not NOT_6193(g23278,g20283);
  not NOT_6194(g23279,g21037);
  not NOT_6195(g23282,g20330);
  not NOT_6196(g23283,g20785);
  not NOT_6197(g23284,g20785);
  not NOT_6198(g23285,g20887);
  not NOT_6199(g23289,g20924);
  not NOT_6200(g23290,g20924);
  not NOT_6201(g23291,g21070);
  not NOT_6202(I22400,g19620);
  not NOT_6203(g23299,I22400);
  not NOT_6204(g23300,g20283);
  not NOT_6205(g23301,g21037);
  not NOT_6206(g23302,g20330);
  not NOT_6207(g23303,g20785);
  not NOT_6208(g23304,g20785);
  not NOT_6209(g23305,g20391);
  not NOT_6210(g23306,g20924);
  not NOT_6211(g23307,g20924);
  not NOT_6212(g23308,g21024);
  not NOT_6213(g23312,g21070);
  not NOT_6214(g23313,g21070);
  not NOT_6215(I22419,g19638);
  not NOT_6216(g23320,I22419);
  not NOT_6217(I22422,g19330);
  not NOT_6218(g23321,I22422);
  not NOT_6219(I22425,g19379);
  not NOT_6220(g23322,I22425);
  not NOT_6221(g23323,g20283);
  not NOT_6222(g23331,g20905);
  not NOT_6223(g23332,g20785);
  not NOT_6224(g23333,g20785);
  not NOT_6225(g23334,g20785);
  not NOT_6226(g23335,g20391);
  not NOT_6227(g23336,g20924);
  not NOT_6228(g23337,g20924);
  not NOT_6229(g23338,g20453);
  not NOT_6230(g23339,g21070);
  not NOT_6231(g23340,g21070);
  not NOT_6232(g23341,g21163);
  not NOT_6233(I22444,g19626);
  not NOT_6234(g23347,I22444);
  not NOT_6235(g23350,g20785);
  not NOT_6236(g23351,g20924);
  not NOT_6237(g23352,g20924);
  not NOT_6238(g23353,g20924);
  not NOT_6239(g23354,g20453);
  not NOT_6240(g23355,g21070);
  not NOT_6241(g23356,g21070);
  not NOT_6242(I22458,g18954);
  not NOT_6243(g23359,I22458);
  not NOT_6244(I22461,g21225);
  not NOT_6245(g23360,I22461);
  not NOT_6246(I22464,g21222);
  not NOT_6247(g23361,I22464);
  not NOT_6248(I22467,g19662);
  not NOT_6249(g23362,I22467);
  not NOT_6250(I22470,g21326);
  not NOT_6251(g23363,I22470);
  not NOT_6252(g23375,g20924);
  not NOT_6253(g23376,g21070);
  not NOT_6254(g23377,g21070);
  not NOT_6255(g23378,g21070);
  not NOT_6256(g23380,g20619);
  not NOT_6257(g23382,g20682);
  not NOT_6258(I22485,g21308);
  not NOT_6259(g23384,I22485);
  not NOT_6260(I22488,g18984);
  not NOT_6261(g23385,I22488);
  not NOT_6262(g23388,g21070);
  not NOT_6263(g23390,g21468);
  not NOT_6264(g23391,g20645);
  not NOT_6265(g23393,g20739);
  not NOT_6266(I22499,g21160);
  not NOT_6267(g23394,I22499);
  not NOT_6268(I22502,g19376);
  not NOT_6269(g23395,I22502);
  not NOT_6270(g23398,g21468);
  not NOT_6271(g23399,g21514);
  not NOT_6272(g23400,g20676);
  not NOT_6273(g23402,g20875);
  not NOT_6274(I22512,g19389);
  not NOT_6275(g23403,I22512);
  not NOT_6276(g23406,g20330);
  not NOT_6277(g23408,g21468);
  not NOT_6278(g23409,g21514);
  not NOT_6279(g23410,g21562);
  not NOT_6280(g23411,g20734);
  not NOT_6281(g23413,g21012);
  not NOT_6282(I22525,g19345);
  not NOT_6283(g23414,I22525);
  not NOT_6284(g23417,g20391);
  not NOT_6285(g23418,g21468);
  not NOT_6286(g23419,g21468);
  not NOT_6287(g23420,g21514);
  not NOT_6288(g23421,g21562);
  not NOT_6289(g23422,g21611);
  not NOT_6290(g23423,g20871);
  not NOT_6291(g23425,g20751);
  not NOT_6292(I22539,g19606);
  not NOT_6293(g23426,I22539);
  not NOT_6294(I22542,g19773);
  not NOT_6295(g23427,I22542);
  not NOT_6296(g23429,g20453);
  not NOT_6297(I22547,g20720);
  not NOT_6298(g23430,I22547);
  not NOT_6299(g23431,g21514);
  not NOT_6300(g23432,g21514);
  not NOT_6301(g23433,g21562);
  not NOT_6302(g23434,g21611);
  not NOT_6303(g23435,g18833);
  not NOT_6304(I22557,g20695);
  not NOT_6305(g23440,I22557);
  not NOT_6306(g23443,g21468);
  not NOT_6307(I22561,g20841);
  not NOT_6308(g23444,I22561);
  not NOT_6309(I22564,g20857);
  not NOT_6310(g23445,I22564);
  not NOT_6311(g23446,g21562);
  not NOT_6312(g23447,g21562);
  not NOT_6313(g23448,g21611);
  not NOT_6314(g23449,g18833);
  not NOT_6315(I22571,g20097);
  not NOT_6316(g23450,I22571);
  not NOT_6317(g23452,g21468);
  not NOT_6318(I22576,g21282);
  not NOT_6319(g23453,I22576);
  not NOT_6320(g23456,g21514);
  not NOT_6321(I22580,g20982);
  not NOT_6322(g23457,I22580);
  not NOT_6323(I22583,g20998);
  not NOT_6324(g23458,I22583);
  not NOT_6325(g23459,g21611);
  not NOT_6326(g23460,g21611);
  not NOT_6327(g23461,g18833);
  not NOT_6328(I22589,g21340);
  not NOT_6329(g23462,I22589);
  not NOT_6330(g23472,g21062);
  not NOT_6331(g23473,g20785);
  not NOT_6332(g23476,g21468);
  not NOT_6333(g23477,g21468);
  not NOT_6334(g23478,g21514);
  not NOT_6335(g23479,g21562);
  not NOT_6336(I22601,g21127);
  not NOT_6337(g23480,I22601);
  not NOT_6338(I22604,g21143);
  not NOT_6339(g23481,I22604);
  not NOT_6340(g23482,g18833);
  not NOT_6341(g23483,g18833);
  not NOT_6342(g23485,g20785);
  not NOT_6343(g23486,g20785);
  not NOT_6344(g23487,g20924);
  not NOT_6345(g23488,g21468);
  not NOT_6346(g23489,g21468);
  not NOT_6347(g23490,g21514);
  not NOT_6348(g23491,g21514);
  not NOT_6349(g23492,g21562);
  not NOT_6350(g23493,g21611);
  not NOT_6351(I22619,g21193);
  not NOT_6352(g23494,I22619);
  not NOT_6353(I22622,g21209);
  not NOT_6354(g23495,I22622);
  not NOT_6355(g23496,g20248);
  not NOT_6356(g23499,g20785);
  not NOT_6357(g23500,g20924);
  not NOT_6358(g23501,g20924);
  not NOT_6359(g23502,g21070);
  not NOT_6360(g23503,g21468);
  not NOT_6361(g23504,g21468);
  not NOT_6362(g23505,g21514);
  not NOT_6363(g23506,g21514);
  not NOT_6364(g23507,g21562);
  not NOT_6365(g23508,g21562);
  not NOT_6366(g23509,g21611);
  not NOT_6367(g23510,g18833);
  not NOT_6368(I22640,g21256);
  not NOT_6369(g23511,I22640);
  not NOT_6370(g23512,g20248);
  not NOT_6371(g23515,g20785);
  not NOT_6372(g23516,g20924);
  not NOT_6373(g23517,g21070);
  not NOT_6374(g23518,g21070);
  not NOT_6375(g23519,g21468);
  not NOT_6376(g23520,g21468);
  not NOT_6377(g23521,g21468);
  not NOT_6378(g23522,g21514);
  not NOT_6379(g23523,g21514);
  not NOT_6380(g23524,g21562);
  not NOT_6381(g23525,g21562);
  not NOT_6382(g23526,g21611);
  not NOT_6383(g23527,g21611);
  not NOT_6384(g23528,g18833);
  not NOT_6385(g23529,g20558);
  not NOT_6386(g23530,g20248);
  not NOT_6387(I22665,g21308);
  not NOT_6388(g23534,I22665);
  not NOT_6389(g23537,g20785);
  not NOT_6390(g23538,g20924);
  not NOT_6391(g23539,g21070);
  not NOT_6392(g23541,g21514);
  not NOT_6393(g23542,g21514);
  not NOT_6394(g23543,g21514);
  not NOT_6395(g23544,g21562);
  not NOT_6396(g23545,g21562);
  not NOT_6397(g23546,g21611);
  not NOT_6398(g23547,g21611);
  not NOT_6399(g23548,g18833);
  not NOT_6400(g23549,g18833);
  not NOT_6401(g23550,g20248);
  not NOT_6402(I22692,g21308);
  not NOT_6403(g23555,I22692);
  not NOT_6404(g23558,g20924);
  not NOT_6405(g23559,g21070);
  not NOT_6406(g23563,g20682);
  not NOT_6407(g23565,g21562);
  not NOT_6408(g23566,g21562);
  not NOT_6409(g23567,g21562);
  not NOT_6410(g23568,g21611);
  not NOT_6411(g23569,g21611);
  not NOT_6412(g23570,g18833);
  not NOT_6413(g23571,g18833);
  not NOT_6414(g23573,g20248);
  not NOT_6415(I22725,g21250);
  not NOT_6416(g23578,I22725);
  not NOT_6417(I22729,g21308);
  not NOT_6418(g23582,I22729);
  not NOT_6419(g23585,g21070);
  not NOT_6420(g23589,g21468);
  not NOT_6421(g23605,g20739);
  not NOT_6422(g23607,g21611);
  not NOT_6423(g23608,g21611);
  not NOT_6424(g23609,g21611);
  not NOT_6425(g23610,g18833);
  not NOT_6426(g23611,g18833);
  not NOT_6427(I22745,g19458);
  not NOT_6428(g23612,I22745);
  not NOT_6429(I22748,g19458);
  not NOT_6430(g23613,I22748);
  not NOT_6431(g23614,g20248);
  not NOT_6432(I22769,g21277);
  not NOT_6433(g23620,I22769);
  not NOT_6434(g23629,g21514);
  not NOT_6435(g23645,g20875);
  not NOT_6436(g23647,g18833);
  not NOT_6437(g23648,g18833);
  not NOT_6438(g23649,g18833);
  not NOT_6439(g23650,g20653);
  not NOT_6440(g23651,g20655);
  not NOT_6441(I22785,g18940);
  not NOT_6442(g23652,I22785);
  not NOT_6443(I22788,g18940);
  not NOT_6444(g23653,I22788);
  not NOT_6445(g23654,g20248);
  not NOT_6446(g23665,g21562);
  not NOT_6447(g23681,g21012);
  not NOT_6448(I22816,g19862);
  not NOT_6449(g23683,I22816);
  not NOT_6450(I22819,g19862);
  not NOT_6451(g23684,I22819);
  not NOT_6452(g23698,g21611);
  not NOT_6453(g23714,g20751);
  not NOT_6454(g23715,g20764);
  not NOT_6455(g23732,g18833);
  not NOT_6456(g23745,g20900);
  not NOT_6457(g23746,g20902);
  not NOT_6458(g23749,g18997);
  not NOT_6459(I22886,g18926);
  not NOT_6460(g23759,I22886);
  not NOT_6461(I22889,g18926);
  not NOT_6462(g23760,I22889);
  not NOT_6463(g23764,g21308);
  not NOT_6464(g23767,g18997);
  not NOT_6465(g23768,g18997);
  not NOT_6466(g23769,g19074);
  not NOT_6467(g23776,g21177);
  not NOT_6468(I22918,g21451);
  not NOT_6469(g23777,I22918);
  not NOT_6470(g23787,g18997);
  not NOT_6471(g23788,g18997);
  not NOT_6472(g23789,g21308);
  not NOT_6473(g23792,g19074);
  not NOT_6474(g23793,g19074);
  not NOT_6475(g23794,g19147);
  not NOT_6476(g23800,g21246);
  not NOT_6477(g23812,g18997);
  not NOT_6478(g23813,g18997);
  not NOT_6479(g23814,g19074);
  not NOT_6480(g23815,g19074);
  not NOT_6481(g23816,g21308);
  not NOT_6482(g23819,g19147);
  not NOT_6483(g23820,g19147);
  not NOT_6484(g23821,g19210);
  not NOT_6485(I22989,g21175);
  not NOT_6486(g23823,I22989);
  not NOT_6487(g23824,g21271);
  not NOT_6488(g23838,g18997);
  not NOT_6489(g23839,g18997);
  not NOT_6490(g23840,g19074);
  not NOT_6491(g23841,g19074);
  not NOT_6492(g23842,g19147);
  not NOT_6493(g23843,g19147);
  not NOT_6494(g23844,g21308);
  not NOT_6495(g23847,g19210);
  not NOT_6496(g23848,g19210);
  not NOT_6497(g23849,g19277);
  not NOT_6498(g23858,g18997);
  not NOT_6499(g23859,g19074);
  not NOT_6500(g23860,g19074);
  not NOT_6501(g23861,g19147);
  not NOT_6502(g23862,g19147);
  not NOT_6503(g23863,g19210);
  not NOT_6504(g23864,g19210);
  not NOT_6505(g23865,g21308);
  not NOT_6506(g23868,g19277);
  not NOT_6507(g23869,g19277);
  not NOT_6508(g23870,g21293);
  not NOT_6509(g23874,g18997);
  not NOT_6510(g23875,g18997);
  not NOT_6511(g23876,g19074);
  not NOT_6512(g23877,g19147);
  not NOT_6513(g23878,g19147);
  not NOT_6514(g23879,g19210);
  not NOT_6515(g23880,g19210);
  not NOT_6516(g23881,g19277);
  not NOT_6517(g23882,g19277);
  not NOT_6518(g23886,g21468);
  not NOT_6519(g23887,g18997);
  not NOT_6520(g23888,g18997);
  not NOT_6521(g23889,g20682);
  not NOT_6522(g23893,g19074);
  not NOT_6523(g23894,g19074);
  not NOT_6524(g23895,g19147);
  not NOT_6525(g23896,g19210);
  not NOT_6526(g23897,g19210);
  not NOT_6527(g23898,g19277);
  not NOT_6528(g23899,g19277);
  not NOT_6529(g23902,g21468);
  not NOT_6530(g23903,g18997);
  not NOT_6531(g23904,g18997);
  not NOT_6532(g23905,g21514);
  not NOT_6533(g23906,g19074);
  not NOT_6534(g23907,g19074);
  not NOT_6535(g23908,g20739);
  not NOT_6536(g23912,g19147);
  not NOT_6537(g23913,g19147);
  not NOT_6538(g23914,g19210);
  not NOT_6539(g23915,g19277);
  not NOT_6540(g23916,g19277);
  not NOT_6541(g23922,g18997);
  not NOT_6542(g23923,g18997);
  not NOT_6543(g23924,g18997);
  not NOT_6544(g23925,g21514);
  not NOT_6545(g23926,g19074);
  not NOT_6546(g23927,g19074);
  not NOT_6547(g23928,g21562);
  not NOT_6548(g23929,g19147);
  not NOT_6549(g23930,g19147);
  not NOT_6550(g23931,g20875);
  not NOT_6551(g23935,g19210);
  not NOT_6552(g23936,g19210);
  not NOT_6553(g23937,g19277);
  not NOT_6554(g23938,g18997);
  not NOT_6555(g23939,g19074);
  not NOT_6556(g23940,g19074);
  not NOT_6557(g23941,g19074);
  not NOT_6558(g23942,g21562);
  not NOT_6559(g23943,g19147);
  not NOT_6560(g23944,g19147);
  not NOT_6561(g23945,g21611);
  not NOT_6562(g23946,g19210);
  not NOT_6563(g23947,g19210);
  not NOT_6564(g23948,g21012);
  not NOT_6565(g23952,g19277);
  not NOT_6566(g23953,g19277);
  not NOT_6567(I23099,g20682);
  not NOT_6568(g23954,I23099);
  not NOT_6569(g23961,g19074);
  not NOT_6570(g23962,g19147);
  not NOT_6571(g23963,g19147);
  not NOT_6572(g23964,g19147);
  not NOT_6573(g23965,g21611);
  not NOT_6574(g23966,g19210);
  not NOT_6575(g23967,g19210);
  not NOT_6576(g23968,g18833);
  not NOT_6577(g23969,g19277);
  not NOT_6578(g23970,g19277);
  not NOT_6579(g23971,g20751);
  not NOT_6580(g23982,g19147);
  not NOT_6581(g23983,g19210);
  not NOT_6582(g23984,g19210);
  not NOT_6583(g23985,g19210);
  not NOT_6584(g23986,g18833);
  not NOT_6585(g23987,g19277);
  not NOT_6586(g23988,g19277);
  not NOT_6587(g23992,g19210);
  not NOT_6588(g23993,g19277);
  not NOT_6589(g23994,g19277);
  not NOT_6590(g23995,g19277);
  not NOT_6591(g23999,g21468);
  not NOT_6592(g24000,g19277);
  not NOT_6593(g24003,g21514);
  not NOT_6594(I23149,g19061);
  not NOT_6595(g24005,I23149);
  not NOT_6596(g24010,g21562);
  not NOT_6597(g24013,g21611);
  not NOT_6598(g24017,g18833);
  not NOT_6599(g24019,g19968);
  not NOT_6600(g24020,g20014);
  not NOT_6601(g24021,g20841);
  not NOT_6602(g24022,g20982);
  not NOT_6603(g24023,g21127);
  not NOT_6604(g24024,g21193);
  not NOT_6605(g24025,g21256);
  not NOT_6606(g24026,g19919);
  not NOT_6607(g24027,g20014);
  not NOT_6608(g24028,g20841);
  not NOT_6609(g24029,g20982);
  not NOT_6610(g24030,g21127);
  not NOT_6611(g24031,g21193);
  not NOT_6612(g24032,g21256);
  not NOT_6613(g24033,g19919);
  not NOT_6614(g24034,g19968);
  not NOT_6615(g24035,g20841);
  not NOT_6616(g24036,g20982);
  not NOT_6617(g24037,g21127);
  not NOT_6618(g24038,g21193);
  not NOT_6619(g24039,g21256);
  not NOT_6620(g24040,g19919);
  not NOT_6621(g24041,g19968);
  not NOT_6622(g24042,g20014);
  not NOT_6623(g24043,g20982);
  not NOT_6624(g24044,g21127);
  not NOT_6625(g24045,g21193);
  not NOT_6626(g24046,g21256);
  not NOT_6627(g24047,g19919);
  not NOT_6628(g24048,g19968);
  not NOT_6629(g24049,g20014);
  not NOT_6630(g24050,g20841);
  not NOT_6631(g24051,g21127);
  not NOT_6632(g24052,g21193);
  not NOT_6633(g24053,g21256);
  not NOT_6634(g24054,g19919);
  not NOT_6635(g24055,g19968);
  not NOT_6636(g24056,g20014);
  not NOT_6637(g24057,g20841);
  not NOT_6638(g24058,g20982);
  not NOT_6639(g24059,g21193);
  not NOT_6640(g24060,g21256);
  not NOT_6641(g24061,g19919);
  not NOT_6642(g24062,g19968);
  not NOT_6643(g24063,g20014);
  not NOT_6644(g24064,g20841);
  not NOT_6645(g24065,g20982);
  not NOT_6646(g24066,g21127);
  not NOT_6647(g24067,g21256);
  not NOT_6648(g24068,g19919);
  not NOT_6649(g24069,g19968);
  not NOT_6650(g24070,g20014);
  not NOT_6651(g24071,g20841);
  not NOT_6652(g24072,g20982);
  not NOT_6653(g24073,g21127);
  not NOT_6654(g24074,g21193);
  not NOT_6655(g24075,g19935);
  not NOT_6656(g24076,g19984);
  not NOT_6657(g24077,g20720);
  not NOT_6658(g24078,g20857);
  not NOT_6659(g24079,g20998);
  not NOT_6660(g24080,g21143);
  not NOT_6661(g24081,g21209);
  not NOT_6662(g24082,g19890);
  not NOT_6663(g24083,g19984);
  not NOT_6664(g24084,g20720);
  not NOT_6665(g24085,g20857);
  not NOT_6666(g24086,g20998);
  not NOT_6667(g24087,g21143);
  not NOT_6668(g24088,g21209);
  not NOT_6669(g24089,g19890);
  not NOT_6670(g24090,g19935);
  not NOT_6671(g24091,g20720);
  not NOT_6672(g24092,g20857);
  not NOT_6673(g24093,g20998);
  not NOT_6674(g24094,g21143);
  not NOT_6675(g24095,g21209);
  not NOT_6676(g24096,g19890);
  not NOT_6677(g24097,g19935);
  not NOT_6678(g24098,g19984);
  not NOT_6679(g24099,g20720);
  not NOT_6680(g24100,g20857);
  not NOT_6681(g24101,g20998);
  not NOT_6682(g24102,g21143);
  not NOT_6683(g24103,g21209);
  not NOT_6684(g24104,g19890);
  not NOT_6685(g24105,g19935);
  not NOT_6686(g24106,g19984);
  not NOT_6687(g24107,g20857);
  not NOT_6688(g24108,g20998);
  not NOT_6689(g24109,g21143);
  not NOT_6690(g24110,g21209);
  not NOT_6691(g24111,g19890);
  not NOT_6692(g24112,g19935);
  not NOT_6693(g24113,g19984);
  not NOT_6694(g24114,g20720);
  not NOT_6695(g24115,g20998);
  not NOT_6696(g24116,g21143);
  not NOT_6697(g24117,g21209);
  not NOT_6698(g24118,g19890);
  not NOT_6699(g24119,g19935);
  not NOT_6700(g24120,g19984);
  not NOT_6701(g24121,g20720);
  not NOT_6702(g24122,g20857);
  not NOT_6703(g24123,g21143);
  not NOT_6704(g24124,g21209);
  not NOT_6705(g24125,g19890);
  not NOT_6706(g24126,g19935);
  not NOT_6707(g24127,g19984);
  not NOT_6708(g24128,g20720);
  not NOT_6709(g24129,g20857);
  not NOT_6710(g24130,g20998);
  not NOT_6711(g24131,g21209);
  not NOT_6712(g24132,g19890);
  not NOT_6713(g24133,g19935);
  not NOT_6714(g24134,g19984);
  not NOT_6715(g24135,g20720);
  not NOT_6716(g24136,g20857);
  not NOT_6717(g24137,g20998);
  not NOT_6718(g24138,g21143);
  not NOT_6719(g24146,g19422);
  not NOT_6720(g24147,g19402);
  not NOT_6721(g24149,g19338);
  not NOT_6722(g24150,g19268);
  not NOT_6723(I23300,g21665);
  not NOT_6724(g24152,I23300);
  not NOT_6725(I23303,g21669);
  not NOT_6726(g24153,I23303);
  not NOT_6727(I23306,g21673);
  not NOT_6728(g24154,I23306);
  not NOT_6729(I23309,g21677);
  not NOT_6730(g24155,I23309);
  not NOT_6731(I23312,g21681);
  not NOT_6732(g24156,I23312);
  not NOT_6733(I23315,g21685);
  not NOT_6734(g24157,I23315);
  not NOT_6735(I23318,g21689);
  not NOT_6736(g24158,I23318);
  not NOT_6737(I23321,g21693);
  not NOT_6738(g24159,I23321);
  not NOT_6739(I23324,g21697);
  not NOT_6740(g24160,I23324);
  not NOT_6741(I23327,g22647);
  not NOT_6742(g24161,I23327);
  not NOT_6743(I23330,g22658);
  not NOT_6744(g24162,I23330);
  not NOT_6745(I23333,g22683);
  not NOT_6746(g24163,I23333);
  not NOT_6747(I23336,g22721);
  not NOT_6748(g24164,I23336);
  not NOT_6749(I23339,g23232);
  not NOT_6750(g24165,I23339);
  not NOT_6751(I23342,g23299);
  not NOT_6752(g24166,I23342);
  not NOT_6753(I23345,g23320);
  not NOT_6754(g24167,I23345);
  not NOT_6755(I23348,g23384);
  not NOT_6756(g24168,I23348);
  not NOT_6757(I23351,g23263);
  not NOT_6758(g24169,I23351);
  not NOT_6759(I23354,g23277);
  not NOT_6760(g24170,I23354);
  not NOT_6761(I23357,g23359);
  not NOT_6762(g24171,I23357);
  not NOT_6763(I23360,g23360);
  not NOT_6764(g24172,I23360);
  not NOT_6765(I23363,g23385);
  not NOT_6766(g24173,I23363);
  not NOT_6767(I23366,g23321);
  not NOT_6768(g24174,I23366);
  not NOT_6769(I23369,g23347);
  not NOT_6770(g24175,I23369);
  not NOT_6771(I23372,g23361);
  not NOT_6772(g24176,I23372);
  not NOT_6773(I23375,g23403);
  not NOT_6774(g24177,I23375);
  not NOT_6775(I23378,g23426);
  not NOT_6776(g24178,I23378);
  not NOT_6777(I23381,g23322);
  not NOT_6778(g24179,I23381);
  not NOT_6779(I23384,g23362);
  not NOT_6780(g24180,I23384);
  not NOT_6781(I23387,g23394);
  not NOT_6782(g24181,I23387);
  not NOT_6783(I23390,g23395);
  not NOT_6784(g24182,I23390);
  not NOT_6785(I23393,g23414);
  not NOT_6786(g24183,I23393);
  not NOT_6787(I23396,g23427);
  not NOT_6788(g24184,I23396);
  not NOT_6789(I23399,g23450);
  not NOT_6790(g24185,I23399);
  not NOT_6791(g24356,g22594);
  not NOT_6792(g24357,g22325);
  not NOT_6793(g24358,g22550);
  not NOT_6794(g24359,g22550);
  not NOT_6795(g24360,g22228);
  not NOT_6796(g24361,g22885);
  not NOT_6797(g24364,g22722);
  not NOT_6798(g24365,g22594);
  not NOT_6799(g24366,g22594);
  not NOT_6800(g24367,g22550);
  not NOT_6801(g24368,g22228);
  not NOT_6802(g24372,g22885);
  not NOT_6803(g24373,g22908);
  not NOT_6804(g24375,g22722);
  not NOT_6805(g24376,g22722);
  not NOT_6806(g24377,g22594);
  not NOT_6807(g24379,g22550);
  not NOT_6808(g24384,g22885);
  not NOT_6809(g24385,g22908);
  not NOT_6810(g24386,g22594);
  not NOT_6811(g24388,g22885);
  not NOT_6812(g24389,g22908);
  not NOT_6813(g24394,g22228);
  not NOT_6814(g24396,g22885);
  not NOT_6815(g24397,g22908);
  not NOT_6816(g24404,g22908);
  not NOT_6817(g24405,g22722);
  not NOT_6818(g24407,g22594);
  not NOT_6819(g24417,g22171);
  not NOT_6820(g24418,g22722);
  not NOT_6821(g24419,g22722);
  not NOT_6822(g24424,g22722);
  not NOT_6823(g24425,g22722);
  not NOT_6824(g24426,g22722);
  not NOT_6825(g24428,g22722);
  not NOT_6826(g24429,g22722);
  not NOT_6827(g24431,g22722);
  not NOT_6828(g24437,g22654);
  not NOT_6829(g24438,g22722);
  not NOT_6830(g24452,g22722);
  not NOT_6831(g24463,g23578);
  not NOT_6832(I23671,g23202);
  not NOT_6833(g24466,I23671);
  not NOT_6834(g24474,g23620);
  not NOT_6835(I23680,g23219);
  not NOT_6836(g24477,I23680);
  not NOT_6837(I23684,g23230);
  not NOT_6838(g24481,I23684);
  not NOT_6839(I23688,g23244);
  not NOT_6840(g24483,I23688);
  not NOT_6841(I23694,g23252);
  not NOT_6842(g24489,I23694);
  not NOT_6843(g24490,g22594);
  not NOT_6844(g24505,g22689);
  not NOT_6845(I23711,g23192);
  not NOT_6846(g24506,I23711);
  not NOT_6847(g24509,g22689);
  not NOT_6848(g24515,g22689);
  not NOT_6849(g24516,g22670);
  not NOT_6850(g24522,g22689);
  not NOT_6851(g24524,g22876);
  not NOT_6852(g24525,g22670);
  not NOT_6853(g24526,g22942);
  not NOT_6854(g24527,g22670);
  not NOT_6855(g24533,g22876);
  not NOT_6856(g24534,g22670);
  not NOT_6857(g24535,g22942);
  not NOT_6858(g24540,g22942);
  not NOT_6859(g24548,g22942);
  not NOT_6860(g24560,g22942);
  not NOT_6861(g24568,g22942);
  not NOT_6862(g24571,g22942);
  not NOT_6863(g24579,g23067);
  not NOT_6864(g24585,g23063);
  not NOT_6865(g24586,g23067);
  not NOT_6866(g24587,g23112);
  not NOT_6867(g24603,g23108);
  not NOT_6868(g24604,g23112);
  not NOT_6869(g24605,g23139);
  not NOT_6870(g24623,g23076);
  not NOT_6871(g24625,g23135);
  not NOT_6872(g24626,g23139);
  not NOT_6873(g24636,g23121);
  not NOT_6874(g24648,g23148);
  not NOT_6875(g24655,g23067);
  not NOT_6876(g24665,g23067);
  not NOT_6877(g24667,g23112);
  not NOT_6878(g24683,g23112);
  not NOT_6879(g24685,g23139);
  not NOT_6880(g24699,g23047);
  not NOT_6881(g24711,g23139);
  not NOT_6882(g24718,g22182);
  not NOT_6883(g24732,g23042);
  not NOT_6884(g24744,g22202);
  not NOT_6885(g24756,g22763);
  not NOT_6886(g24759,g23003);
  not NOT_6887(g24770,g22763);
  not NOT_6888(g24778,g23286);
  not NOT_6889(g24789,g23309);
  not NOT_6890(g24791,g23850);
  not NOT_6891(g24795,g23342);
  not NOT_6892(g24818,g23191);
  not NOT_6893(I23998,g22182);
  not NOT_6894(g24819,I23998);
  not NOT_6895(g24825,g23204);
  not NOT_6896(I24008,g22182);
  not NOT_6897(g24836,I24008);
  not NOT_6898(g24839,g23436);
  not NOT_6899(I24022,g22182);
  not NOT_6900(g24850,I24022);
  not NOT_6901(I24038,g22202);
  not NOT_6902(g24866,I24038);
  not NOT_6903(I24041,g22182);
  not NOT_6904(g24869,I24041);
  not NOT_6905(g24891,g23231);
  not NOT_6906(I24060,g22202);
  not NOT_6907(g24893,I24060);
  not NOT_6908(I24078,g22360);
  not NOT_6909(g24911,I24078);
  not NOT_6910(I24089,g22409);
  not NOT_6911(g24920,I24089);
  not NOT_6912(g24960,g23716);
  not NOT_6913(g24963,g22342);
  not NOT_6914(I24128,g23009);
  not NOT_6915(g24964,I24128);
  not NOT_6916(g24966,g22763);
  not NOT_6917(g24971,g23590);
  not NOT_6918(g24978,g22342);
  not NOT_6919(g24979,g22369);
  not NOT_6920(g24980,g22384);
  not NOT_6921(g24981,g22763);
  not NOT_6922(g24982,g22763);
  not NOT_6923(g24985,g23586);
  not NOT_6924(g24986,g23590);
  not NOT_6925(g24987,g23630);
  not NOT_6926(g24991,g22369);
  not NOT_6927(g24992,g22417);
  not NOT_6928(g24993,g22384);
  not NOT_6929(g24994,g22432);
  not NOT_6930(g24995,g22763);
  not NOT_6931(g24996,g22763);
  not NOT_6932(g24999,g23626);
  not NOT_6933(g25000,g23630);
  not NOT_6934(g25001,g23666);
  not NOT_6935(g25006,g22417);
  not NOT_6936(g25007,g22457);
  not NOT_6937(g25008,g22432);
  not NOT_6938(g25009,g22472);
  not NOT_6939(g25011,g22763);
  not NOT_6940(g25013,g23599);
  not NOT_6941(g25015,g23662);
  not NOT_6942(g25016,g23666);
  not NOT_6943(g25017,g23699);
  not NOT_6944(g25023,g22457);
  not NOT_6945(g25024,g22472);
  not NOT_6946(g25025,g22498);
  not NOT_6947(I24191,g22360);
  not NOT_6948(g25027,I24191);
  not NOT_6949(g25032,g23639);
  not NOT_6950(g25034,g23695);
  not NOT_6951(g25035,g23699);
  not NOT_6952(g25036,g23733);
  not NOT_6953(g25039,g22498);
  not NOT_6954(g25044,g23675);
  not NOT_6955(g25046,g23729);
  not NOT_6956(g25047,g23733);
  not NOT_6957(I24215,g22360);
  not NOT_6958(g25051,I24215);
  not NOT_6959(g25055,g23590);
  not NOT_6960(g25060,g23708);
  not NOT_6961(I24228,g22409);
  not NOT_6962(g25064,I24228);
  not NOT_6963(g25070,g23590);
  not NOT_6964(g25072,g23630);
  not NOT_6965(I24237,g23823);
  not NOT_6966(g25073,I24237);
  not NOT_6967(g25080,g23742);
  not NOT_6968(g25081,g22342);
  not NOT_6969(g25082,g22342);
  not NOT_6970(g25083,g23782);
  not NOT_6971(g25090,g23630);
  not NOT_6972(g25092,g23666);
  not NOT_6973(g25097,g22342);
  not NOT_6974(g25098,g22369);
  not NOT_6975(g25099,g22369);
  not NOT_6976(g25100,g22384);
  not NOT_6977(g25101,g22384);
  not NOT_6978(g25109,g23666);
  not NOT_6979(g25111,g23699);
  not NOT_6980(I24278,g23440);
  not NOT_6981(g25114,I24278);
  not NOT_6982(I24281,g23440);
  not NOT_6983(g25115,I24281);
  not NOT_6984(g25116,g22369);
  not NOT_6985(g25117,g22417);
  not NOT_6986(g25118,g22417);
  not NOT_6987(g25119,g22384);
  not NOT_6988(g25120,g22432);
  not NOT_6989(g25121,g22432);
  not NOT_6990(g25131,g23699);
  not NOT_6991(g25133,g23733);
  not NOT_6992(g25134,g22417);
  not NOT_6993(g25135,g22457);
  not NOT_6994(g25136,g22457);
  not NOT_6995(g25137,g22432);
  not NOT_6996(g25138,g22472);
  not NOT_6997(g25139,g22472);
  not NOT_6998(g25140,g22228);
  not NOT_6999(g25153,g23733);
  not NOT_7000(g25154,g22457);
  not NOT_7001(g25155,g22472);
  not NOT_7002(g25156,g22498);
  not NOT_7003(g25157,g22498);
  not NOT_7004(g25158,g22228);
  not NOT_7005(I24331,g22976);
  not NOT_7006(g25167,I24331);
  not NOT_7007(I24334,g22976);
  not NOT_7008(g25168,I24334);
  not NOT_7009(g25169,g22763);
  not NOT_7010(g25170,g22498);
  not NOT_7011(g25171,g22228);
  not NOT_7012(g25174,g23890);
  not NOT_7013(g25180,g23529);
  not NOT_7014(g25182,g22763);
  not NOT_7015(g25183,g22763);
  not NOT_7016(g25184,g22763);
  not NOT_7017(g25185,g22228);
  not NOT_7018(g25188,g23909);
  not NOT_7019(g25193,g22763);
  not NOT_7020(g25194,g22763);
  not NOT_7021(g25195,g22763);
  not NOT_7022(g25196,g22763);
  not NOT_7023(g25197,g23958);
  not NOT_7024(g25198,g22228);
  not NOT_7025(g25202,g23932);
  not NOT_7026(g25206,g23613);
  not NOT_7027(g25208,g22763);
  not NOT_7028(g25209,g22763);
  not NOT_7029(g25210,g23802);
  not NOT_7030(g25211,g22763);
  not NOT_7031(g25212,g22763);
  not NOT_7032(g25213,g23293);
  not NOT_7033(g25214,g22228);
  not NOT_7034(g25218,g23949);
  not NOT_7035(I24393,g23453);
  not NOT_7036(g25219,I24393);
  not NOT_7037(I24396,g23453);
  not NOT_7038(g25220,I24396);
  not NOT_7039(g25221,g23653);
  not NOT_7040(I24400,g23954);
  not NOT_7041(g25222,I24400);
  not NOT_7042(g25224,g22763);
  not NOT_7043(g25225,g23802);
  not NOT_7044(g25226,g22763);
  not NOT_7045(g25227,g22763);
  not NOT_7046(g25228,g23828);
  not NOT_7047(g25230,g23314);
  not NOT_7048(g25231,g22228);
  not NOT_7049(g25232,g22228);
  not NOT_7050(g25239,g23972);
  not NOT_7051(g25240,g23650);
  not NOT_7052(g25241,g23651);
  not NOT_7053(g25242,g23684);
  not NOT_7054(g25243,g22763);
  not NOT_7055(g25244,g23802);
  not NOT_7056(g25245,g22763);
  not NOT_7057(g25246,g23828);
  not NOT_7058(g25248,g22228);
  not NOT_7059(g25249,g22228);
  not NOT_7060(I24434,g22763);
  not NOT_7061(g25250,I24434);
  not NOT_7062(I24445,g22923);
  not NOT_7063(g25259,I24445);
  not NOT_7064(I24448,g22923);
  not NOT_7065(g25260,I24448);
  not NOT_7066(g25262,g22763);
  not NOT_7067(g25263,g22763);
  not NOT_7068(g25264,g23828);
  not NOT_7069(I24455,g22541);
  not NOT_7070(g25265,I24455);
  not NOT_7071(g25266,g22228);
  not NOT_7072(g25267,g22228);
  not NOT_7073(g25272,g23715);
  not NOT_7074(g25273,g23978);
  not NOT_7075(g25274,g22763);
  not NOT_7076(g25282,g22763);
  not NOT_7077(g25283,g22763);
  not NOT_7078(I24474,g22546);
  not NOT_7079(g25284,I24474);
  not NOT_7080(g25286,g22228);
  not NOT_7081(g25287,g22228);
  not NOT_7082(g25288,g22228);
  not NOT_7083(g25289,g22228);
  not NOT_7084(g25296,g23745);
  not NOT_7085(g25297,g23746);
  not NOT_7086(g25298,g23760);
  not NOT_7087(g25299,g22763);
  not NOT_7088(g25307,g22763);
  not NOT_7089(g25308,g22763);
  not NOT_7090(g25316,g22763);
  not NOT_7091(I24497,g22592);
  not NOT_7092(g25322,I24497);
  not NOT_7093(g25324,g22228);
  not NOT_7094(g25325,g22228);
  not NOT_7095(g25326,g22228);
  not NOT_7096(g25327,g22161);
  not NOT_7097(g25340,g22763);
  not NOT_7098(g25348,g22763);
  not NOT_7099(g25356,g22763);
  not NOT_7100(g25369,g22228);
  not NOT_7101(g25370,g22228);
  not NOT_7102(g25380,g23776);
  not NOT_7103(g25388,g22763);
  not NOT_7104(g25399,g22763);
  not NOT_7105(g25409,g22228);
  not NOT_7106(g25410,g22228);
  not NOT_7107(I24558,g23777);
  not NOT_7108(g25423,I24558);
  not NOT_7109(g25424,g23800);
  not NOT_7110(g25438,g22763);
  not NOT_7111(g25451,g22228);
  not NOT_7112(g25452,g22228);
  not NOT_7113(g25465,g23824);
  not NOT_7114(g25480,g22228);
  not NOT_7115(g25481,g22228);
  not NOT_7116(g25505,g22228);
  not NOT_7117(g25506,g22228);
  not NOT_7118(g25513,g23870);
  not NOT_7119(g25517,g22228);
  not NOT_7120(g25523,g22550);
  not NOT_7121(g25524,g22228);
  not NOT_7122(g25525,g22550);
  not NOT_7123(g25528,g22594);
  not NOT_7124(g25529,g22763);
  not NOT_7125(g25533,g22550);
  not NOT_7126(g25534,g22763);
  not NOT_7127(g25535,g22763);
  not NOT_7128(g25538,g22594);
  not NOT_7129(g25541,g22763);
  not NOT_7130(g25542,g22763);
  not NOT_7131(g25544,g22594);
  not NOT_7132(g25546,g22550);
  not NOT_7133(g25547,g22550);
  not NOT_7134(g25548,g22550);
  not NOT_7135(g25549,g22763);
  not NOT_7136(g25550,g22763);
  not NOT_7137(g25552,g22594);
  not NOT_7138(g25553,g22550);
  not NOT_7139(g25554,g22550);
  not NOT_7140(g25555,g22550);
  not NOT_7141(g25556,g22763);
  not NOT_7142(g25557,g22763);
  not NOT_7143(g25558,g22594);
  not NOT_7144(g25560,g22550);
  not NOT_7145(g25561,g22550);
  not NOT_7146(g25562,g22763);
  not NOT_7147(g25563,g22594);
  not NOT_7148(g25564,g22312);
  not NOT_7149(g25566,g22550);
  not NOT_7150(I24759,g24229);
  not NOT_7151(g25620,I24759);
  not NOT_7152(I24781,g24264);
  not NOT_7153(g25640,I24781);
  not NOT_7154(I24784,g24265);
  not NOT_7155(g25641,I24784);
  not NOT_7156(I24787,g24266);
  not NOT_7157(g25642,I24787);
  not NOT_7158(I24839,g24298);
  not NOT_7159(g25692,I24839);
  not NOT_7160(g25766,g24439);
  not NOT_7161(I24920,g25513);
  not NOT_7162(g25771,I24920);
  not NOT_7163(g25773,g24453);
  not NOT_7164(g25781,g24510);
  not NOT_7165(g25783,g25250);
  not NOT_7166(g25786,g24518);
  not NOT_7167(g25790,g25027);
  not NOT_7168(g25820,g25051);
  not NOT_7169(g25830,g24485);
  not NOT_7170(g25837,g25064);
  not NOT_7171(g25838,g25250);
  not NOT_7172(g25849,g24491);
  not NOT_7173(g25869,g25250);
  not NOT_7174(g25882,g25026);
  not NOT_7175(g25886,g24537);
  not NOT_7176(g25892,g24528);
  not NOT_7177(g25893,g24541);
  not NOT_7178(g25899,g24997);
  not NOT_7179(I25005,g24417);
  not NOT_7180(g25903,I25005);
  not NOT_7181(I25028,g24484);
  not NOT_7182(g25930,I25028);
  not NOT_7183(g25994,g24575);
  not NOT_7184(I25095,g25265);
  not NOT_7185(g25997,I25095);
  not NOT_7186(I25105,g25284);
  not NOT_7187(g26026,I25105);
  not NOT_7188(g26054,g24804);
  not NOT_7189(I25115,g25322);
  not NOT_7190(g26055,I25115);
  not NOT_7191(g26081,g24619);
  not NOT_7192(g26083,g24809);
  not NOT_7193(g26093,g24814);
  not NOT_7194(I25146,g24911);
  not NOT_7195(g26105,I25146);
  not NOT_7196(I25161,g24920);
  not NOT_7197(g26131,I25161);
  not NOT_7198(I25190,g25423);
  not NOT_7199(g26187,I25190);
  not NOT_7200(g26260,g24759);
  not NOT_7201(g26284,g24875);
  not NOT_7202(g26326,g24872);
  not NOT_7203(g26337,g24818);
  not NOT_7204(g26340,g24953);
  not NOT_7205(I25327,g24641);
  not NOT_7206(g26364,I25327);
  not NOT_7207(I25351,g24466);
  not NOT_7208(g26400,I25351);
  not NOT_7209(I25356,g24374);
  not NOT_7210(g26424,I25356);
  not NOT_7211(I25359,g24715);
  not NOT_7212(g26483,I25359);
  not NOT_7213(I25366,g24477);
  not NOT_7214(g26488,I25366);
  not NOT_7215(I25369,g24891);
  not NOT_7216(g26510,I25369);
  not NOT_7217(g26518,g25233);
  not NOT_7218(I25380,g24481);
  not NOT_7219(g26519,I25380);
  not NOT_7220(g26548,g25255);
  not NOT_7221(I25391,g24483);
  not NOT_7222(g26549,I25391);
  not NOT_7223(g26575,g25268);
  not NOT_7224(I25399,g24489);
  not NOT_7225(g26576,I25399);
  not NOT_7226(g26605,g25293);
  not NOT_7227(g26607,g25382);
  not NOT_7228(g26608,g25334);
  not NOT_7229(g26614,g25426);
  not NOT_7230(g26615,g25432);
  not NOT_7231(g26631,g25467);
  not NOT_7232(g26632,g25473);
  not NOT_7233(g26634,g25317);
  not NOT_7234(g26648,g25115);
  not NOT_7235(g26653,g25337);
  not NOT_7236(g26654,g25275);
  not NOT_7237(g26655,g25492);
  not NOT_7238(g26656,g25495);
  not NOT_7239(g26672,g25275);
  not NOT_7240(g26679,g25385);
  not NOT_7241(g26680,g25300);
  not NOT_7242(g26681,g25396);
  not NOT_7243(g26682,g25309);
  not NOT_7244(g26683,g25514);
  not NOT_7245(g26693,g25300);
  not NOT_7246(g26700,g25429);
  not NOT_7247(g26701,g25341);
  not NOT_7248(g26702,g25309);
  not NOT_7249(g26709,g25435);
  not NOT_7250(g26710,g25349);
  not NOT_7251(g26718,g25168);
  not NOT_7252(g26720,g25275);
  not NOT_7253(g26724,g25341);
  not NOT_7254(g26731,g25470);
  not NOT_7255(g26732,g25389);
  not NOT_7256(g26736,g25349);
  not NOT_7257(g26743,g25476);
  not NOT_7258(g26744,g25400);
  not NOT_7259(g26754,g25300);
  not NOT_7260(g26758,g25389);
  not NOT_7261(g26765,g25309);
  not NOT_7262(g26769,g25400);
  not NOT_7263(g26776,g25498);
  not NOT_7264(g26777,g25439);
  not NOT_7265(g26784,g25341);
  not NOT_7266(g26788,g25349);
  not NOT_7267(g26792,g25439);
  not NOT_7268(I25511,g25073);
  not NOT_7269(g26801,I25511);
  not NOT_7270(I25514,g25073);
  not NOT_7271(g26802,I25514);
  not NOT_7272(g26803,g25389);
  not NOT_7273(g26804,g25400);
  not NOT_7274(g26810,g25220);
  not NOT_7275(g26811,g25206);
  not NOT_7276(g26812,g25439);
  not NOT_7277(g26814,g25221);
  not NOT_7278(g26816,g25260);
  not NOT_7279(g26817,g25242);
  not NOT_7280(I25530,g25222);
  not NOT_7281(g26818,I25530);
  not NOT_7282(I25534,g25448);
  not NOT_7283(g26820,I25534);
  not NOT_7284(g26824,g25298);
  not NOT_7285(I25541,g25180);
  not NOT_7286(g26825,I25541);
  not NOT_7287(g26827,g24819);
  not NOT_7288(g26830,g24411);
  not NOT_7289(g26831,g24836);
  not NOT_7290(g26832,g24850);
  not NOT_7291(I25552,g25240);
  not NOT_7292(g26834,I25552);
  not NOT_7293(I25555,g25241);
  not NOT_7294(g26835,I25555);
  not NOT_7295(g26836,g24866);
  not NOT_7296(g26837,g24869);
  not NOT_7297(I25562,g25250);
  not NOT_7298(g26840,I25562);
  not NOT_7299(g26841,g24893);
  not NOT_7300(I25567,g25272);
  not NOT_7301(g26843,I25567);
  not NOT_7302(I25576,g25296);
  not NOT_7303(g26850,I25576);
  not NOT_7304(I25579,g25297);
  not NOT_7305(g26851,I25579);
  not NOT_7306(I25586,g25537);
  not NOT_7307(g26856,I25586);
  not NOT_7308(I25591,g25380);
  not NOT_7309(g26859,I25591);
  not NOT_7310(I25594,g25531);
  not NOT_7311(g26860,I25594);
  not NOT_7312(I25598,g25424);
  not NOT_7313(g26862,I25598);
  not NOT_7314(g26869,g24842);
  not NOT_7315(I25606,g25465);
  not NOT_7316(g26870,I25606);
  not NOT_7317(I25677,g25640);
  not NOT_7318(g26935,I25677);
  not NOT_7319(I25680,g25641);
  not NOT_7320(g26936,I25680);
  not NOT_7321(I25683,g25642);
  not NOT_7322(g26937,I25683);
  not NOT_7323(I25689,g25688);
  not NOT_7324(g26941,I25689);
  not NOT_7325(I25692,g25689);
  not NOT_7326(g26942,I25692);
  not NOT_7327(I25695,g25690);
  not NOT_7328(g26943,I25695);
  not NOT_7329(g26973,g26105);
  not NOT_7330(g26987,g26131);
  not NOT_7331(g26990,g26105);
  not NOT_7332(g27004,g26131);
  not NOT_7333(g27009,g25911);
  not NOT_7334(g27011,g25917);
  not NOT_7335(I25743,g25903);
  not NOT_7336(g27013,I25743);
  not NOT_7337(g27014,g25888);
  not NOT_7338(g27015,g26869);
  not NOT_7339(g27017,g25895);
  not NOT_7340(I25750,g26823);
  not NOT_7341(g27018,I25750);
  not NOT_7342(g27038,g25932);
  not NOT_7343(I25779,g26424);
  not NOT_7344(g27051,I25779);
  not NOT_7345(I25786,g26424);
  not NOT_7346(g27064,I25786);
  not NOT_7347(I25790,g26424);
  not NOT_7348(g27074,I25790);
  not NOT_7349(g27084,g26673);
  not NOT_7350(g27088,g26694);
  not NOT_7351(g27089,g26703);
  not NOT_7352(g27091,g26725);
  not NOT_7353(g27092,g26737);
  not NOT_7354(g27100,g26759);
  not NOT_7355(g27101,g26770);
  not NOT_7356(g27112,g26793);
  not NOT_7357(g27142,g26105);
  not NOT_7358(g27155,g26131);
  not NOT_7359(I25869,g25851);
  not NOT_7360(g27163,I25869);
  not NOT_7361(I25882,g25776);
  not NOT_7362(g27187,I25882);
  not NOT_7363(g27237,g26162);
  not NOT_7364(g27242,g26183);
  not NOT_7365(g27245,g26209);
  not NOT_7366(g27279,g26330);
  not NOT_7367(I26004,g26818);
  not NOT_7368(g27320,I26004);
  not NOT_7369(g27349,g26352);
  not NOT_7370(I26100,g26365);
  not NOT_7371(g27402,I26100);
  not NOT_7372(g27415,g26382);
  not NOT_7373(I26130,g26510);
  not NOT_7374(g27438,I26130);
  not NOT_7375(g27492,g26598);
  not NOT_7376(I26195,g26260);
  not NOT_7377(g27527,I26195);
  not NOT_7378(g27554,g26625);
  not NOT_7379(g27565,g26645);
  not NOT_7380(g27573,g26667);
  not NOT_7381(g27576,g26081);
  not NOT_7382(g27583,g26686);
  not NOT_7383(g27585,g25994);
  not NOT_7384(g27592,g26715);
  not NOT_7385(g27597,g26745);
  not NOT_7386(I26296,g26820);
  not NOT_7387(g27662,I26296);
  not NOT_7388(I26309,g26825);
  not NOT_7389(g27675,I26309);
  not NOT_7390(g27698,g26648);
  not NOT_7391(I26334,g26834);
  not NOT_7392(g27708,I26334);
  not NOT_7393(I26337,g26835);
  not NOT_7394(g27709,I26337);
  not NOT_7395(g27730,g26424);
  not NOT_7396(I26356,g26843);
  not NOT_7397(g27736,I26356);
  not NOT_7398(g27737,g26718);
  not NOT_7399(I26378,g26850);
  not NOT_7400(g27773,I26378);
  not NOT_7401(I26381,g26851);
  not NOT_7402(g27774,I26381);
  not NOT_7403(g27830,g26802);
  not NOT_7404(I26406,g26187);
  not NOT_7405(g27831,I26406);
  not NOT_7406(I26409,g26187);
  not NOT_7407(g27832,I26409);
  not NOT_7408(I26427,g26859);
  not NOT_7409(g27880,I26427);
  not NOT_7410(I26430,g26856);
  not NOT_7411(g27881,I26430);
  not NOT_7412(g27928,g26810);
  not NOT_7413(I26448,g26860);
  not NOT_7414(g27929,I26448);
  not NOT_7415(I26451,g26862);
  not NOT_7416(g27930,I26451);
  not NOT_7417(I26466,g26870);
  not NOT_7418(g27956,I26466);
  not NOT_7419(g27961,g26816);
  not NOT_7420(I26479,g25771);
  not NOT_7421(g27967,I26479);
  not NOT_7422(g27971,g26673);
  not NOT_7423(g27975,g26694);
  not NOT_7424(g27976,g26703);
  not NOT_7425(g27977,g26105);
  not NOT_7426(g27983,g26725);
  not NOT_7427(g27984,g26737);
  not NOT_7428(g27985,g26131);
  not NOT_7429(g27989,g26759);
  not NOT_7430(g27990,g26770);
  not NOT_7431(g27991,g25852);
  not NOT_7432(I26503,g26811);
  not NOT_7433(g27993,I26503);
  not NOT_7434(g27994,g26793);
  not NOT_7435(I26508,g26814);
  not NOT_7436(g27996,I26508);
  not NOT_7437(I26512,g26817);
  not NOT_7438(g27998,I26512);
  not NOT_7439(I26516,g26824);
  not NOT_7440(g28009,I26516);
  not NOT_7441(g28032,g26365);
  not NOT_7442(g28033,g26365);
  not NOT_7443(g28034,g26365);
  not NOT_7444(g28036,g26365);
  not NOT_7445(g28037,g26365);
  not NOT_7446(g28038,g26365);
  not NOT_7447(g28039,g26365);
  not NOT_7448(g28040,g26365);
  not NOT_7449(I26578,g26941);
  not NOT_7450(g28079,I26578);
  not NOT_7451(I26581,g26942);
  not NOT_7452(g28080,I26581);
  not NOT_7453(I26584,g26943);
  not NOT_7454(g28081,I26584);
  not NOT_7455(g28119,g27008);
  not NOT_7456(g28120,g27108);
  not NOT_7457(g28121,g27093);
  not NOT_7458(g28126,g27122);
  not NOT_7459(g28127,g27102);
  not NOT_7460(I26638,g27965);
  not NOT_7461(g28137,I26638);
  not NOT_7462(I26649,g27675);
  not NOT_7463(g28142,I26649);
  not NOT_7464(I26654,g27576);
  not NOT_7465(g28147,I26654);
  not NOT_7466(I26664,g27708);
  not NOT_7467(g28155,I26664);
  not NOT_7468(I26667,g27585);
  not NOT_7469(g28156,I26667);
  not NOT_7470(I26670,g27709);
  not NOT_7471(g28157,I26670);
  not NOT_7472(I26676,g27736);
  not NOT_7473(g28161,I26676);
  not NOT_7474(I26679,g27773);
  not NOT_7475(g28162,I26679);
  not NOT_7476(I26682,g27774);
  not NOT_7477(g28163,I26682);
  not NOT_7478(I26687,g27880);
  not NOT_7479(g28166,I26687);
  not NOT_7480(I26693,g27930);
  not NOT_7481(g28173,I26693);
  not NOT_7482(I26700,g27956);
  not NOT_7483(g28181,I26700);
  not NOT_7484(I26705,g27967);
  not NOT_7485(g28184,I26705);
  not NOT_7486(I26710,g27511);
  not NOT_7487(g28187,I26710);
  not NOT_7488(g28241,g27064);
  not NOT_7489(g28250,g27074);
  not NOT_7490(I26785,g27013);
  not NOT_7491(g28262,I26785);
  not NOT_7492(I26799,g27660);
  not NOT_7493(g28274,I26799);
  not NOT_7494(g28294,g27295);
  not NOT_7495(g28307,g27306);
  not NOT_7496(g28321,g27317);
  not NOT_7497(g28325,g27463);
  not NOT_7498(g28326,g27414);
  not NOT_7499(I26880,g27527);
  not NOT_7500(g28367,I26880);
  not NOT_7501(g28370,g27528);
  not NOT_7502(g28380,g27064);
  not NOT_7503(g28399,g27074);
  not NOT_7504(I26925,g27015);
  not NOT_7505(g28431,I26925);
  not NOT_7506(I26929,g27980);
  not NOT_7507(g28436,I26929);
  not NOT_7508(g28441,g27629);
  not NOT_7509(I26936,g27599);
  not NOT_7510(g28443,I26936);
  not NOT_7511(I26952,g27972);
  not NOT_7512(g28463,I26952);
  not NOT_7513(g28479,g27654);
  not NOT_7514(I26989,g27277);
  not NOT_7515(g28508,I26989);
  not NOT_7516(g28559,g27700);
  not NOT_7517(g28575,g27711);
  not NOT_7518(g28579,g27714);
  not NOT_7519(g28590,g27724);
  not NOT_7520(g28593,g27727);
  not NOT_7521(g28598,g27717);
  not NOT_7522(g28604,g27759);
  not NOT_7523(g28606,g27762);
  not NOT_7524(g28608,g27670);
  not NOT_7525(g28615,g27817);
  not NOT_7526(g28620,g27679);
  not NOT_7527(g28633,g27687);
  not NOT_7528(g28648,g27693);
  not NOT_7529(g28656,g27742);
  not NOT_7530(g28669,g27705);
  not NOT_7531(g28675,g27779);
  not NOT_7532(g28678,g27800);
  not NOT_7533(g28693,g27837);
  not NOT_7534(g28696,g27858);
  not NOT_7535(I27192,g27662);
  not NOT_7536(g28709,I27192);
  not NOT_7537(g28711,g27886);
  not NOT_7538(g28713,g27907);
  not NOT_7539(g28726,g27937);
  not NOT_7540(I27232,g27993);
  not NOT_7541(g28752,I27232);
  not NOT_7542(I27235,g27320);
  not NOT_7543(g28753,I27235);
  not NOT_7544(I27238,g27320);
  not NOT_7545(g28754,I27238);
  not NOT_7546(I27253,g27996);
  not NOT_7547(g28779,I27253);
  not NOT_7548(I27271,g27998);
  not NOT_7549(g28819,I27271);
  not NOT_7550(I27314,g28009);
  not NOT_7551(g28917,I27314);
  not NOT_7552(g28918,g27832);
  not NOT_7553(g28954,g27830);
  not NOT_7554(I27368,g27881);
  not NOT_7555(g29013,I27368);
  not NOT_7556(g29014,g27742);
  not NOT_7557(I27385,g27438);
  not NOT_7558(g29041,I27385);
  not NOT_7559(I27388,g27698);
  not NOT_7560(g29042,I27388);
  not NOT_7561(I27391,g27929);
  not NOT_7562(g29043,I27391);
  not NOT_7563(g29044,g27742);
  not NOT_7564(g29045,g27779);
  not NOT_7565(g29056,g27800);
  not NOT_7566(I27401,g27051);
  not NOT_7567(g29067,I27401);
  not NOT_7568(g29079,g27742);
  not NOT_7569(g29080,g27779);
  not NOT_7570(g29081,g27837);
  not NOT_7571(g29092,g27800);
  not NOT_7572(g29093,g27858);
  not NOT_7573(g29115,g27779);
  not NOT_7574(g29116,g27837);
  not NOT_7575(g29117,g27886);
  not NOT_7576(g29128,g27800);
  not NOT_7577(g29129,g27858);
  not NOT_7578(g29130,g27907);
  not NOT_7579(I27449,g27737);
  not NOT_7580(g29147,I27449);
  not NOT_7581(g29149,g27837);
  not NOT_7582(g29150,g27886);
  not NOT_7583(g29151,g27858);
  not NOT_7584(g29152,g27907);
  not NOT_7585(g29153,g27937);
  not NOT_7586(g29169,g27886);
  not NOT_7587(g29170,g27907);
  not NOT_7588(g29171,g27937);
  not NOT_7589(g29172,g27020);
  not NOT_7590(g29177,g27937);
  not NOT_7591(I27481,g27928);
  not NOT_7592(g29185,I27481);
  not NOT_7593(g29190,g27046);
  not NOT_7594(I27492,g27511);
  not NOT_7595(g29194,I27492);
  not NOT_7596(I27495,g27961);
  not NOT_7597(g29195,I27495);
  not NOT_7598(g29196,g27059);
  not NOT_7599(I27543,g28187);
  not NOT_7600(g29209,I27543);
  not NOT_7601(I27546,g29041);
  not NOT_7602(g29210,I27546);
  not NOT_7603(I27549,g28161);
  not NOT_7604(g29211,I27549);
  not NOT_7605(I27552,g28162);
  not NOT_7606(g29212,I27552);
  not NOT_7607(I27555,g28142);
  not NOT_7608(g29213,I27555);
  not NOT_7609(I27558,g28155);
  not NOT_7610(g29214,I27558);
  not NOT_7611(I27561,g28163);
  not NOT_7612(g29215,I27561);
  not NOT_7613(I27564,g28166);
  not NOT_7614(g29216,I27564);
  not NOT_7615(I27567,g28181);
  not NOT_7616(g29217,I27567);
  not NOT_7617(I27570,g28262);
  not NOT_7618(g29218,I27570);
  not NOT_7619(I27573,g28157);
  not NOT_7620(g29219,I27573);
  not NOT_7621(I27576,g28173);
  not NOT_7622(g29220,I27576);
  not NOT_7623(I27579,g28184);
  not NOT_7624(g29221,I27579);
  not NOT_7625(g29310,g28991);
  not NOT_7626(g29311,g28998);
  not NOT_7627(g29312,g28877);
  not NOT_7628(I27677,g28156);
  not NOT_7629(g29317,I27677);
  not NOT_7630(g29318,g29029);
  not NOT_7631(g29333,g28167);
  not NOT_7632(g29339,g28274);
  not NOT_7633(g29342,g28188);
  not NOT_7634(g29343,g28174);
  not NOT_7635(g29348,g28194);
  not NOT_7636(I27713,g28224);
  not NOT_7637(g29353,I27713);
  not NOT_7638(I27718,g28231);
  not NOT_7639(g29358,I27718);
  not NOT_7640(g29365,g29067);
  not NOT_7641(I27730,g28752);
  not NOT_7642(g29368,I27730);
  not NOT_7643(I27735,g28779);
  not NOT_7644(g29371,I27735);
  not NOT_7645(I27738,g28140);
  not NOT_7646(g29372,I27738);
  not NOT_7647(I27742,g28819);
  not NOT_7648(g29374,I27742);
  not NOT_7649(I27749,g28917);
  not NOT_7650(g29379,I27749);
  not NOT_7651(g29385,g28180);
  not NOT_7652(I27758,g28119);
  not NOT_7653(g29474,I27758);
  not NOT_7654(I27777,g29043);
  not NOT_7655(g29491,I27777);
  not NOT_7656(I27784,g29013);
  not NOT_7657(g29498,I27784);
  not NOT_7658(g29505,g29186);
  not NOT_7659(g29507,g28353);
  not NOT_7660(g29597,g28444);
  not NOT_7661(I27927,g28803);
  not NOT_7662(g29653,I27927);
  not NOT_7663(I27941,g28803);
  not NOT_7664(g29669,I27941);
  not NOT_7665(I27954,g28803);
  not NOT_7666(g29689,I27954);
  not NOT_7667(g29697,g28336);
  not NOT_7668(g29707,g28504);
  not NOT_7669(I27970,g28803);
  not NOT_7670(g29713,I27970);
  not NOT_7671(g29725,g28349);
  not NOT_7672(g29744,g28431);
  not NOT_7673(g29745,g28500);
  not NOT_7674(I28002,g28153);
  not NOT_7675(g29755,I28002);
  not NOT_7676(I28014,g28158);
  not NOT_7677(g29765,I28014);
  not NOT_7678(g29800,g28363);
  not NOT_7679(g29811,g28376);
  not NOT_7680(g29812,g28381);
  not NOT_7681(I28062,g29194);
  not NOT_7682(g29814,I28062);
  not NOT_7683(g29846,g28391);
  not NOT_7684(g29847,g28395);
  not NOT_7685(g29862,g28406);
  not NOT_7686(g29863,g28410);
  not NOT_7687(g29878,g28421);
  not NOT_7688(g29893,g28755);
  not NOT_7689(I28128,g28314);
  not NOT_7690(g29897,I28128);
  not NOT_7691(g29905,g28783);
  not NOT_7692(g29906,g28793);
  not NOT_7693(g29911,g28780);
  not NOT_7694(g29912,g28827);
  not NOT_7695(g29913,g28840);
  not NOT_7696(g29920,g28824);
  not NOT_7697(g29921,g28864);
  not NOT_7698(g29922,g28837);
  not NOT_7699(g29923,g28874);
  not NOT_7700(g29925,g28820);
  not NOT_7701(g29927,g28861);
  not NOT_7702(g29928,g28871);
  not NOT_7703(g29929,g28914);
  not NOT_7704(I28162,g28803);
  not NOT_7705(g29930,I28162);
  not NOT_7706(g29939,g28857);
  not NOT_7707(g29941,g28900);
  not NOT_7708(g29942,g28867);
  not NOT_7709(g29944,g28911);
  not NOT_7710(I28174,g28803);
  not NOT_7711(g29945,I28174);
  not NOT_7712(g29948,g28853);
  not NOT_7713(g29950,g28896);
  not NOT_7714(g29953,g28907);
  not NOT_7715(g29955,g28950);
  not NOT_7716(I28185,g28803);
  not NOT_7717(g29956,I28185);
  not NOT_7718(g29960,g28885);
  not NOT_7719(g29961,g28892);
  not NOT_7720(g29963,g28931);
  not NOT_7721(g29965,g28903);
  not NOT_7722(g29967,g28946);
  not NOT_7723(I28199,g28803);
  not NOT_7724(g29970,I28199);
  not NOT_7725(g29976,g29018);
  not NOT_7726(g29977,g28920);
  not NOT_7727(g29978,g28927);
  not NOT_7728(g29980,g28935);
  not NOT_7729(g29981,g28942);
  not NOT_7730(g29983,g28977);
  not NOT_7731(g29993,g29018);
  not NOT_7732(g29994,g29049);
  not NOT_7733(g29995,g28955);
  not NOT_7734(g29996,g28962);
  not NOT_7735(g29997,g29060);
  not NOT_7736(g29998,g28966);
  not NOT_7737(g29999,g28973);
  not NOT_7738(I28241,g28709);
  not NOT_7739(g30012,I28241);
  not NOT_7740(g30016,g29049);
  not NOT_7741(g30017,g29085);
  not NOT_7742(g30018,g28987);
  not NOT_7743(g30019,g29060);
  not NOT_7744(g30020,g29097);
  not NOT_7745(g30021,g28994);
  not NOT_7746(g30022,g29001);
  not NOT_7747(g30036,g29085);
  not NOT_7748(g30037,g29121);
  not NOT_7749(g30038,g29097);
  not NOT_7750(g30039,g29134);
  not NOT_7751(g30040,g29025);
  not NOT_7752(g30052,g29018);
  not NOT_7753(g30053,g29121);
  not NOT_7754(g30054,g29134);
  not NOT_7755(g30055,g29157);
  not NOT_7756(g30063,g29015);
  not NOT_7757(g30065,g29049);
  not NOT_7758(g30067,g29060);
  not NOT_7759(g30068,g29157);
  not NOT_7760(I28301,g29042);
  not NOT_7761(g30072,I28301);
  not NOT_7762(g30074,g29046);
  not NOT_7763(g30076,g29085);
  not NOT_7764(g30077,g29057);
  not NOT_7765(g30079,g29097);
  not NOT_7766(g30085,g29082);
  not NOT_7767(g30087,g29121);
  not NOT_7768(g30088,g29094);
  not NOT_7769(g30090,g29134);
  not NOT_7770(g30097,g29118);
  not NOT_7771(g30100,g29131);
  not NOT_7772(g30102,g29157);
  not NOT_7773(I28336,g29147);
  not NOT_7774(g30105,I28336);
  not NOT_7775(g30113,g29154);
  not NOT_7776(I28349,g28367);
  not NOT_7777(g30116,I28349);
  not NOT_7778(g30142,g28754);
  not NOT_7779(I28390,g29185);
  not NOT_7780(g30155,I28390);
  not NOT_7781(I28419,g29195);
  not NOT_7782(g30182,I28419);
  not NOT_7783(g30184,g28144);
  not NOT_7784(I28434,g28114);
  not NOT_7785(g30195,I28434);
  not NOT_7786(g30206,g28436);
  not NOT_7787(I28458,g28443);
  not NOT_7788(g30217,I28458);
  not NOT_7789(g30218,g28918);
  not NOT_7790(I28480,g28652);
  not NOT_7791(g30237,I28480);
  not NOT_7792(g30259,g28463);
  not NOT_7793(g30292,g28736);
  not NOT_7794(I28540,g28954);
  not NOT_7795(g30295,I28540);
  not NOT_7796(g30296,g28889);
  not NOT_7797(g30297,g28758);
  not NOT_7798(g30299,g28765);
  not NOT_7799(I28548,g28147);
  not NOT_7800(g30301,I28548);
  not NOT_7801(g30302,g28924);
  not NOT_7802(g30303,g28786);
  not NOT_7803(g30305,g28939);
  not NOT_7804(g30306,g28796);
  not NOT_7805(g30309,g28959);
  not NOT_7806(g30310,g28830);
  not NOT_7807(g30312,g28970);
  not NOT_7808(g30313,g28843);
  not NOT_7809(g30318,g28274);
  not NOT_7810(I28572,g28274);
  not NOT_7811(g30321,I28572);
  not NOT_7812(g30322,g28431);
  not NOT_7813(I28576,g28431);
  not NOT_7814(g30325,I28576);
  not NOT_7815(I28579,g29474);
  not NOT_7816(g30326,I28579);
  not NOT_7817(I28582,g30116);
  not NOT_7818(g30327,I28582);
  not NOT_7819(I28585,g30217);
  not NOT_7820(g30328,I28585);
  not NOT_7821(I28588,g29368);
  not NOT_7822(g30329,I28588);
  not NOT_7823(I28591,g29371);
  not NOT_7824(g30330,I28591);
  not NOT_7825(I28594,g29379);
  not NOT_7826(g30331,I28594);
  not NOT_7827(I28597,g29374);
  not NOT_7828(g30332,I28597);
  not NOT_7829(I28832,g30301);
  not NOT_7830(g30565,I28832);
  not NOT_7831(g30567,g29930);
  not NOT_7832(g30568,g29339);
  not NOT_7833(I28838,g29372);
  not NOT_7834(g30569,I28838);
  not NOT_7835(g30572,g29945);
  not NOT_7836(g30578,g29956);
  not NOT_7837(I28851,g29317);
  not NOT_7838(g30591,I28851);
  not NOT_7839(g30593,g29970);
  not NOT_7840(I28866,g29730);
  not NOT_7841(g30606,I28866);
  not NOT_7842(I28872,g30072);
  not NOT_7843(g30610,I28872);
  not NOT_7844(I28883,g30105);
  not NOT_7845(g30729,I28883);
  not NOT_7846(I28897,g30155);
  not NOT_7847(g30917,I28897);
  not NOT_7848(I28908,g30182);
  not NOT_7849(g30928,I28908);
  not NOT_7850(I28913,g30322);
  not NOT_7851(g30931,I28913);
  not NOT_7852(g30983,g29657);
  not NOT_7853(g30989,g29672);
  not NOT_7854(g30990,g29676);
  not NOT_7855(I28925,g29987);
  not NOT_7856(g30991,I28925);
  not NOT_7857(g30996,g29694);
  not NOT_7858(g30997,g29702);
  not NOT_7859(g30998,g29719);
  not NOT_7860(g30999,g29722);
  not NOT_7861(g31000,g29737);
  not NOT_7862(g31013,g29679);
  not NOT_7863(g31138,g29778);
  not NOT_7864(I29002,g29675);
  not NOT_7865(g31189,I29002);
  not NOT_7866(I29013,g29705);
  not NOT_7867(g31213,I29013);
  not NOT_7868(g31227,g29744);
  not NOT_7869(g31239,g29916);
  not NOT_7870(g31243,g29933);
  not NOT_7871(I29139,g29382);
  not NOT_7872(g31479,I29139);
  not NOT_7873(I29149,g29384);
  not NOT_7874(g31487,I29149);
  not NOT_7875(I29182,g30012);
  not NOT_7876(g31521,I29182);
  not NOT_7877(I29185,g30012);
  not NOT_7878(g31522,I29185);
  not NOT_7879(I29199,g30237);
  not NOT_7880(g31578,I29199);
  not NOT_7881(I29204,g29505);
  not NOT_7882(g31596,I29204);
  not NOT_7883(I29207,g30293);
  not NOT_7884(g31601,I29207);
  not NOT_7885(g31608,g29653);
  not NOT_7886(I29211,g30298);
  not NOT_7887(g31609,I29211);
  not NOT_7888(I29214,g30300);
  not NOT_7889(g31616,I29214);
  not NOT_7890(g31623,g29669);
  not NOT_7891(I29218,g30304);
  not NOT_7892(g31624,I29218);
  not NOT_7893(I29221,g30307);
  not NOT_7894(g31631,I29221);
  not NOT_7895(g31638,g29689);
  not NOT_7896(I29225,g30311);
  not NOT_7897(g31639,I29225);
  not NOT_7898(I29228,g30314);
  not NOT_7899(g31646,I29228);
  not NOT_7900(g31653,g29713);
  not NOT_7901(I29233,g30295);
  not NOT_7902(g31655,I29233);
  not NOT_7903(I29236,g29498);
  not NOT_7904(g31656,I29236);
  not NOT_7905(I29239,g29498);
  not NOT_7906(g31657,I29239);
  not NOT_7907(I29242,g29313);
  not NOT_7908(g31658,I29242);
  not NOT_7909(I29245,g29491);
  not NOT_7910(g31665,I29245);
  not NOT_7911(I29248,g29491);
  not NOT_7912(g31666,I29248);
  not NOT_7913(g31667,g30142);
  not NOT_7914(I29337,g30286);
  not NOT_7915(g31771,I29337);
  not NOT_7916(I29363,g30218);
  not NOT_7917(g31791,I29363);
  not NOT_7918(I29368,g30321);
  not NOT_7919(g31794,I29368);
  not NOT_7920(I29371,g30325);
  not NOT_7921(g31795,I29371);
  not NOT_7922(g31796,g29385);
  not NOT_7923(g31797,g29385);
  not NOT_7924(g31798,g29385);
  not NOT_7925(g31799,g29385);
  not NOT_7926(g31800,g29385);
  not NOT_7927(g31801,g29385);
  not NOT_7928(g31802,g29385);
  not NOT_7929(g31803,g29385);
  not NOT_7930(g31804,g29385);
  not NOT_7931(g31805,g29385);
  not NOT_7932(g31806,g29385);
  not NOT_7933(g31807,g29385);
  not NOT_7934(g31808,g29385);
  not NOT_7935(g31809,g29385);
  not NOT_7936(g31810,g29385);
  not NOT_7937(g31811,g29385);
  not NOT_7938(g31812,g29385);
  not NOT_7939(g31813,g29385);
  not NOT_7940(g31814,g29385);
  not NOT_7941(g31815,g29385);
  not NOT_7942(g31816,g29385);
  not NOT_7943(g31817,g29385);
  not NOT_7944(g31818,g29385);
  not NOT_7945(g31819,g29385);
  not NOT_7946(g31820,g29385);
  not NOT_7947(g31821,g29385);
  not NOT_7948(g31822,g29385);
  not NOT_7949(g31823,g29385);
  not NOT_7950(g31824,g29385);
  not NOT_7951(g31825,g29385);
  not NOT_7952(g31826,g29385);
  not NOT_7953(g31827,g29385);
  not NOT_7954(g31828,g29385);
  not NOT_7955(g31829,g29385);
  not NOT_7956(g31830,g29385);
  not NOT_7957(g31831,g29385);
  not NOT_7958(g31832,g29385);
  not NOT_7959(g31833,g29385);
  not NOT_7960(g31834,g29385);
  not NOT_7961(g31835,g29385);
  not NOT_7962(g31836,g29385);
  not NOT_7963(g31837,g29385);
  not NOT_7964(g31838,g29385);
  not NOT_7965(g31839,g29385);
  not NOT_7966(g31840,g29385);
  not NOT_7967(g31841,g29385);
  not NOT_7968(g31842,g29385);
  not NOT_7969(g31843,g29385);
  not NOT_7970(g31844,g29385);
  not NOT_7971(g31845,g29385);
  not NOT_7972(g31846,g29385);
  not NOT_7973(g31847,g29385);
  not NOT_7974(g31848,g29385);
  not NOT_7975(g31849,g29385);
  not NOT_7976(g31850,g29385);
  not NOT_7977(g31851,g29385);
  not NOT_7978(g31852,g29385);
  not NOT_7979(g31853,g29385);
  not NOT_7980(g31854,g29385);
  not NOT_7981(g31855,g29385);
  not NOT_7982(g31856,g29385);
  not NOT_7983(g31857,g29385);
  not NOT_7984(g31858,g29385);
  not NOT_7985(g31859,g29385);
  not NOT_7986(I29438,g30610);
  not NOT_7987(g31860,I29438);
  not NOT_7988(I29441,g30917);
  not NOT_7989(g31861,I29441);
  not NOT_7990(I29444,g30928);
  not NOT_7991(g31862,I29444);
  not NOT_7992(I29447,g30729);
  not NOT_7993(g31863,I29447);
  not NOT_7994(g31937,g30991);
  not NOT_7995(g31945,g31189);
  not NOT_7996(I29571,g31783);
  not NOT_7997(g32015,I29571);
  not NOT_7998(I29579,g30565);
  not NOT_7999(g32021,I29579);
  not NOT_8000(I29582,g30591);
  not NOT_8001(g32024,I29582);
  not NOT_8002(I29585,g31655);
  not NOT_8003(g32027,I29585);
  not NOT_8004(g32033,g30929);
  not NOT_8005(g32038,g30934);
  not NOT_8006(g32090,g31003);
  not NOT_8007(g32099,g31009);
  not NOT_8008(g32118,g31008);
  not NOT_8009(g32137,g31134);
  not NOT_8010(g32138,g31233);
  not NOT_8011(I29717,g30931);
  not NOT_8012(g32185,I29717);
  not NOT_8013(I29720,g30931);
  not NOT_8014(g32186,I29720);
  not NOT_8015(g32192,g31262);
  not NOT_8016(g32201,g31509);
  not NOT_8017(g32318,g31596);
  not NOT_8018(g32329,g31522);
  not NOT_8019(I29891,g31578);
  not NOT_8020(g32363,I29891);
  not NOT_8021(I29894,g31771);
  not NOT_8022(g32364,I29894);
  not NOT_8023(g32377,g30984);
  not NOT_8024(I29909,g31791);
  not NOT_8025(g32381,I29909);
  not NOT_8026(g32382,g31657);
  not NOT_8027(I29913,g30605);
  not NOT_8028(g32383,I29913);
  not NOT_8029(g32384,g31666);
  not NOT_8030(g32393,g30922);
  not NOT_8031(g32394,g30601);
  not NOT_8032(I29936,g30606);
  not NOT_8033(g32404,I29936);
  not NOT_8034(I29939,g31667);
  not NOT_8035(g32407,I29939);
  not NOT_8036(g32415,g31591);
  not NOT_8037(g32421,g31213);
  not NOT_8038(g32430,g30984);
  not NOT_8039(I29961,g30984);
  not NOT_8040(g32433,I29961);
  not NOT_8041(g32434,g31189);
  not NOT_8042(I29965,g31189);
  not NOT_8043(g32437,I29965);
  not NOT_8044(g32438,g30991);
  not NOT_8045(I29969,g30991);
  not NOT_8046(g32441,I29969);
  not NOT_8047(g32442,g31213);
  not NOT_8048(I29973,g31213);
  not NOT_8049(g32445,I29973);
  not NOT_8050(g32446,g31596);
  not NOT_8051(I29977,g31596);
  not NOT_8052(g32449,I29977);
  not NOT_8053(g32450,g31591);
  not NOT_8054(I29981,g31591);
  not NOT_8055(g32453,I29981);
  not NOT_8056(g32456,g31376);
  not NOT_8057(g32457,g30735);
  not NOT_8058(g32458,g30825);
  not NOT_8059(g32459,g31070);
  not NOT_8060(g32460,g31194);
  not NOT_8061(g32461,g30614);
  not NOT_8062(g32462,g30673);
  not NOT_8063(g32463,g31566);
  not NOT_8064(g32464,g30735);
  not NOT_8065(g32465,g30825);
  not NOT_8066(g32466,g31070);
  not NOT_8067(g32467,g31194);
  not NOT_8068(g32468,g30614);
  not NOT_8069(g32469,g30673);
  not NOT_8070(g32470,g31566);
  not NOT_8071(g32471,g31376);
  not NOT_8072(g32472,g30825);
  not NOT_8073(g32473,g31070);
  not NOT_8074(g32474,g31194);
  not NOT_8075(g32475,g30614);
  not NOT_8076(g32476,g30673);
  not NOT_8077(g32477,g31566);
  not NOT_8078(g32478,g31376);
  not NOT_8079(g32479,g30735);
  not NOT_8080(g32480,g31070);
  not NOT_8081(g32481,g31194);
  not NOT_8082(g32482,g30614);
  not NOT_8083(g32483,g30673);
  not NOT_8084(g32484,g31566);
  not NOT_8085(g32485,g31376);
  not NOT_8086(g32486,g30735);
  not NOT_8087(g32487,g30825);
  not NOT_8088(g32488,g31194);
  not NOT_8089(g32489,g30614);
  not NOT_8090(g32490,g30673);
  not NOT_8091(g32491,g31566);
  not NOT_8092(g32492,g31376);
  not NOT_8093(g32493,g30735);
  not NOT_8094(g32494,g30825);
  not NOT_8095(g32495,g31070);
  not NOT_8096(g32496,g30614);
  not NOT_8097(g32497,g30673);
  not NOT_8098(g32498,g31566);
  not NOT_8099(g32499,g31376);
  not NOT_8100(g32500,g30735);
  not NOT_8101(g32501,g30825);
  not NOT_8102(g32502,g31070);
  not NOT_8103(g32503,g31194);
  not NOT_8104(g32504,g30673);
  not NOT_8105(g32505,g31566);
  not NOT_8106(g32506,g31376);
  not NOT_8107(g32507,g30735);
  not NOT_8108(g32508,g30825);
  not NOT_8109(g32509,g31070);
  not NOT_8110(g32510,g31194);
  not NOT_8111(g32511,g30614);
  not NOT_8112(g32512,g31566);
  not NOT_8113(g32513,g31376);
  not NOT_8114(g32514,g30735);
  not NOT_8115(g32515,g30825);
  not NOT_8116(g32516,g31070);
  not NOT_8117(g32517,g31194);
  not NOT_8118(g32518,g30614);
  not NOT_8119(g32519,g30673);
  not NOT_8120(g32521,g31376);
  not NOT_8121(g32522,g30735);
  not NOT_8122(g32523,g30825);
  not NOT_8123(g32524,g31070);
  not NOT_8124(g32525,g31170);
  not NOT_8125(g32526,g30614);
  not NOT_8126(g32527,g30673);
  not NOT_8127(g32528,g31554);
  not NOT_8128(g32529,g30735);
  not NOT_8129(g32530,g30825);
  not NOT_8130(g32531,g31070);
  not NOT_8131(g32532,g31170);
  not NOT_8132(g32533,g30614);
  not NOT_8133(g32534,g30673);
  not NOT_8134(g32535,g31554);
  not NOT_8135(g32536,g31376);
  not NOT_8136(g32537,g30825);
  not NOT_8137(g32538,g31070);
  not NOT_8138(g32539,g31170);
  not NOT_8139(g32540,g30614);
  not NOT_8140(g32541,g30673);
  not NOT_8141(g32542,g31554);
  not NOT_8142(g32543,g31376);
  not NOT_8143(g32544,g30735);
  not NOT_8144(g32545,g31070);
  not NOT_8145(g32546,g31170);
  not NOT_8146(g32547,g30614);
  not NOT_8147(g32548,g30673);
  not NOT_8148(g32549,g31554);
  not NOT_8149(g32550,g31376);
  not NOT_8150(g32551,g30735);
  not NOT_8151(g32552,g30825);
  not NOT_8152(g32553,g31170);
  not NOT_8153(g32554,g30614);
  not NOT_8154(g32555,g30673);
  not NOT_8155(g32556,g31554);
  not NOT_8156(g32557,g31376);
  not NOT_8157(g32558,g30735);
  not NOT_8158(g32559,g30825);
  not NOT_8159(g32560,g31070);
  not NOT_8160(g32561,g30614);
  not NOT_8161(g32562,g30673);
  not NOT_8162(g32563,g31554);
  not NOT_8163(g32564,g31376);
  not NOT_8164(g32565,g30735);
  not NOT_8165(g32566,g30825);
  not NOT_8166(g32567,g31070);
  not NOT_8167(g32568,g31170);
  not NOT_8168(g32569,g30673);
  not NOT_8169(g32570,g31554);
  not NOT_8170(g32571,g31376);
  not NOT_8171(g32572,g30735);
  not NOT_8172(g32573,g30825);
  not NOT_8173(g32574,g31070);
  not NOT_8174(g32575,g31170);
  not NOT_8175(g32576,g30614);
  not NOT_8176(g32577,g31554);
  not NOT_8177(g32578,g31376);
  not NOT_8178(g32579,g30735);
  not NOT_8179(g32580,g30825);
  not NOT_8180(g32581,g31070);
  not NOT_8181(g32582,g31170);
  not NOT_8182(g32583,g30614);
  not NOT_8183(g32584,g30673);
  not NOT_8184(g32586,g31376);
  not NOT_8185(g32587,g30735);
  not NOT_8186(g32588,g30825);
  not NOT_8187(g32589,g31070);
  not NOT_8188(g32590,g31154);
  not NOT_8189(g32591,g30614);
  not NOT_8190(g32592,g30673);
  not NOT_8191(g32593,g31542);
  not NOT_8192(g32594,g30735);
  not NOT_8193(g32595,g30825);
  not NOT_8194(g32596,g31070);
  not NOT_8195(g32597,g31154);
  not NOT_8196(g32598,g30614);
  not NOT_8197(g32599,g30673);
  not NOT_8198(g32600,g31542);
  not NOT_8199(g32601,g31376);
  not NOT_8200(g32602,g30825);
  not NOT_8201(g32603,g31070);
  not NOT_8202(g32604,g31154);
  not NOT_8203(g32605,g30614);
  not NOT_8204(g32606,g30673);
  not NOT_8205(g32607,g31542);
  not NOT_8206(g32608,g31376);
  not NOT_8207(g32609,g30735);
  not NOT_8208(g32610,g31070);
  not NOT_8209(g32611,g31154);
  not NOT_8210(g32612,g30614);
  not NOT_8211(g32613,g30673);
  not NOT_8212(g32614,g31542);
  not NOT_8213(g32615,g31376);
  not NOT_8214(g32616,g30735);
  not NOT_8215(g32617,g30825);
  not NOT_8216(g32618,g31154);
  not NOT_8217(g32619,g30614);
  not NOT_8218(g32620,g30673);
  not NOT_8219(g32621,g31542);
  not NOT_8220(g32622,g31376);
  not NOT_8221(g32623,g30735);
  not NOT_8222(g32624,g30825);
  not NOT_8223(g32625,g31070);
  not NOT_8224(g32626,g30614);
  not NOT_8225(g32627,g30673);
  not NOT_8226(g32628,g31542);
  not NOT_8227(g32629,g31376);
  not NOT_8228(g32630,g30735);
  not NOT_8229(g32631,g30825);
  not NOT_8230(g32632,g31070);
  not NOT_8231(g32633,g31154);
  not NOT_8232(g32634,g30673);
  not NOT_8233(g32635,g31542);
  not NOT_8234(g32636,g31376);
  not NOT_8235(g32637,g30735);
  not NOT_8236(g32638,g30825);
  not NOT_8237(g32639,g31070);
  not NOT_8238(g32640,g31154);
  not NOT_8239(g32641,g30614);
  not NOT_8240(g32642,g31542);
  not NOT_8241(g32643,g31376);
  not NOT_8242(g32644,g30735);
  not NOT_8243(g32645,g30825);
  not NOT_8244(g32646,g31070);
  not NOT_8245(g32647,g31154);
  not NOT_8246(g32648,g30614);
  not NOT_8247(g32649,g30673);
  not NOT_8248(g32651,g31376);
  not NOT_8249(g32652,g30735);
  not NOT_8250(g32653,g30825);
  not NOT_8251(g32654,g31070);
  not NOT_8252(g32655,g30614);
  not NOT_8253(g32656,g30673);
  not NOT_8254(g32657,g31528);
  not NOT_8255(g32658,g31579);
  not NOT_8256(g32659,g30735);
  not NOT_8257(g32660,g30825);
  not NOT_8258(g32661,g31070);
  not NOT_8259(g32662,g30614);
  not NOT_8260(g32663,g30673);
  not NOT_8261(g32664,g31528);
  not NOT_8262(g32665,g31579);
  not NOT_8263(g32666,g31376);
  not NOT_8264(g32667,g30825);
  not NOT_8265(g32668,g31070);
  not NOT_8266(g32669,g30614);
  not NOT_8267(g32670,g30673);
  not NOT_8268(g32671,g31528);
  not NOT_8269(g32672,g31579);
  not NOT_8270(g32673,g31376);
  not NOT_8271(g32674,g30735);
  not NOT_8272(g32675,g31070);
  not NOT_8273(g32676,g30614);
  not NOT_8274(g32677,g30673);
  not NOT_8275(g32678,g31528);
  not NOT_8276(g32679,g31579);
  not NOT_8277(g32680,g31376);
  not NOT_8278(g32681,g30735);
  not NOT_8279(g32682,g30825);
  not NOT_8280(g32683,g30614);
  not NOT_8281(g32684,g30673);
  not NOT_8282(g32685,g31528);
  not NOT_8283(g32686,g31579);
  not NOT_8284(g32687,g31376);
  not NOT_8285(g32688,g30735);
  not NOT_8286(g32689,g30825);
  not NOT_8287(g32690,g31070);
  not NOT_8288(g32691,g30673);
  not NOT_8289(g32692,g31528);
  not NOT_8290(g32693,g31579);
  not NOT_8291(g32694,g31376);
  not NOT_8292(g32695,g30735);
  not NOT_8293(g32696,g30825);
  not NOT_8294(g32697,g31070);
  not NOT_8295(g32698,g30614);
  not NOT_8296(g32699,g31528);
  not NOT_8297(g32700,g31579);
  not NOT_8298(g32701,g31376);
  not NOT_8299(g32702,g30735);
  not NOT_8300(g32703,g30825);
  not NOT_8301(g32704,g31070);
  not NOT_8302(g32705,g30614);
  not NOT_8303(g32706,g30673);
  not NOT_8304(g32707,g31579);
  not NOT_8305(g32708,g31376);
  not NOT_8306(g32709,g30735);
  not NOT_8307(g32710,g30825);
  not NOT_8308(g32711,g31070);
  not NOT_8309(g32712,g30614);
  not NOT_8310(g32713,g30673);
  not NOT_8311(g32714,g31528);
  not NOT_8312(g32716,g31376);
  not NOT_8313(g32717,g30735);
  not NOT_8314(g32718,g30825);
  not NOT_8315(g32719,g31672);
  not NOT_8316(g32720,g31710);
  not NOT_8317(g32721,g31021);
  not NOT_8318(g32722,g30937);
  not NOT_8319(g32723,g31327);
  not NOT_8320(g32724,g30735);
  not NOT_8321(g32725,g30825);
  not NOT_8322(g32726,g31672);
  not NOT_8323(g32727,g31710);
  not NOT_8324(g32728,g31021);
  not NOT_8325(g32729,g30937);
  not NOT_8326(g32730,g31327);
  not NOT_8327(g32731,g31376);
  not NOT_8328(g32732,g30825);
  not NOT_8329(g32733,g31672);
  not NOT_8330(g32734,g31710);
  not NOT_8331(g32735,g31021);
  not NOT_8332(g32736,g30937);
  not NOT_8333(g32737,g31327);
  not NOT_8334(g32738,g31376);
  not NOT_8335(g32739,g30735);
  not NOT_8336(g32740,g31672);
  not NOT_8337(g32741,g31710);
  not NOT_8338(g32742,g31021);
  not NOT_8339(g32743,g30937);
  not NOT_8340(g32744,g31327);
  not NOT_8341(g32745,g31376);
  not NOT_8342(g32746,g30735);
  not NOT_8343(g32747,g30825);
  not NOT_8344(g32748,g31710);
  not NOT_8345(g32749,g31021);
  not NOT_8346(g32750,g30937);
  not NOT_8347(g32751,g31327);
  not NOT_8348(g32752,g31376);
  not NOT_8349(g32753,g30735);
  not NOT_8350(g32754,g30825);
  not NOT_8351(g32755,g31672);
  not NOT_8352(g32756,g31021);
  not NOT_8353(g32757,g30937);
  not NOT_8354(g32758,g31327);
  not NOT_8355(g32759,g31376);
  not NOT_8356(g32760,g30735);
  not NOT_8357(g32761,g30825);
  not NOT_8358(g32762,g31672);
  not NOT_8359(g32763,g31710);
  not NOT_8360(g32764,g30937);
  not NOT_8361(g32765,g31327);
  not NOT_8362(g32766,g31376);
  not NOT_8363(g32767,g30735);
  not NOT_8364(g32768,g30825);
  not NOT_8365(g32769,g31672);
  not NOT_8366(g32770,g31710);
  not NOT_8367(g32771,g31021);
  not NOT_8368(g32772,g31327);
  not NOT_8369(g32773,g31376);
  not NOT_8370(g32774,g30735);
  not NOT_8371(g32775,g30825);
  not NOT_8372(g32776,g31672);
  not NOT_8373(g32777,g31710);
  not NOT_8374(g32778,g31021);
  not NOT_8375(g32779,g30937);
  not NOT_8376(g32781,g31376);
  not NOT_8377(g32782,g30735);
  not NOT_8378(g32783,g30825);
  not NOT_8379(g32784,g31672);
  not NOT_8380(g32785,g31710);
  not NOT_8381(g32786,g31021);
  not NOT_8382(g32787,g30937);
  not NOT_8383(g32788,g31327);
  not NOT_8384(g32789,g30735);
  not NOT_8385(g32790,g30825);
  not NOT_8386(g32791,g31672);
  not NOT_8387(g32792,g31710);
  not NOT_8388(g32793,g31021);
  not NOT_8389(g32794,g30937);
  not NOT_8390(g32795,g31327);
  not NOT_8391(g32796,g31376);
  not NOT_8392(g32797,g30825);
  not NOT_8393(g32798,g31672);
  not NOT_8394(g32799,g31710);
  not NOT_8395(g32800,g31021);
  not NOT_8396(g32801,g30937);
  not NOT_8397(g32802,g31327);
  not NOT_8398(g32803,g31376);
  not NOT_8399(g32804,g30735);
  not NOT_8400(g32805,g31672);
  not NOT_8401(g32806,g31710);
  not NOT_8402(g32807,g31021);
  not NOT_8403(g32808,g30937);
  not NOT_8404(g32809,g31327);
  not NOT_8405(g32810,g31376);
  not NOT_8406(g32811,g30735);
  not NOT_8407(g32812,g30825);
  not NOT_8408(g32813,g31710);
  not NOT_8409(g32814,g31021);
  not NOT_8410(g32815,g30937);
  not NOT_8411(g32816,g31327);
  not NOT_8412(g32817,g31376);
  not NOT_8413(g32818,g30735);
  not NOT_8414(g32819,g30825);
  not NOT_8415(g32820,g31672);
  not NOT_8416(g32821,g31021);
  not NOT_8417(g32822,g30937);
  not NOT_8418(g32823,g31327);
  not NOT_8419(g32824,g31376);
  not NOT_8420(g32825,g30735);
  not NOT_8421(g32826,g30825);
  not NOT_8422(g32827,g31672);
  not NOT_8423(g32828,g31710);
  not NOT_8424(g32829,g30937);
  not NOT_8425(g32830,g31327);
  not NOT_8426(g32831,g31376);
  not NOT_8427(g32832,g30735);
  not NOT_8428(g32833,g30825);
  not NOT_8429(g32834,g31672);
  not NOT_8430(g32835,g31710);
  not NOT_8431(g32836,g31021);
  not NOT_8432(g32837,g31327);
  not NOT_8433(g32838,g31376);
  not NOT_8434(g32839,g30735);
  not NOT_8435(g32840,g30825);
  not NOT_8436(g32841,g31672);
  not NOT_8437(g32842,g31710);
  not NOT_8438(g32843,g31021);
  not NOT_8439(g32844,g30937);
  not NOT_8440(g32846,g31376);
  not NOT_8441(g32847,g30735);
  not NOT_8442(g32848,g30825);
  not NOT_8443(g32849,g31021);
  not NOT_8444(g32850,g30937);
  not NOT_8445(g32851,g31327);
  not NOT_8446(g32852,g30614);
  not NOT_8447(g32853,g30673);
  not NOT_8448(g32854,g30735);
  not NOT_8449(g32855,g30825);
  not NOT_8450(g32856,g31021);
  not NOT_8451(g32857,g30937);
  not NOT_8452(g32858,g31327);
  not NOT_8453(g32859,g30614);
  not NOT_8454(g32860,g30673);
  not NOT_8455(g32861,g31376);
  not NOT_8456(g32862,g30825);
  not NOT_8457(g32863,g31021);
  not NOT_8458(g32864,g30937);
  not NOT_8459(g32865,g31327);
  not NOT_8460(g32866,g30614);
  not NOT_8461(g32867,g30673);
  not NOT_8462(g32868,g31376);
  not NOT_8463(g32869,g30735);
  not NOT_8464(g32870,g31021);
  not NOT_8465(g32871,g30937);
  not NOT_8466(g32872,g31327);
  not NOT_8467(g32873,g30614);
  not NOT_8468(g32874,g30673);
  not NOT_8469(g32875,g31376);
  not NOT_8470(g32876,g30735);
  not NOT_8471(g32877,g30825);
  not NOT_8472(g32878,g30937);
  not NOT_8473(g32879,g31327);
  not NOT_8474(g32880,g30614);
  not NOT_8475(g32881,g30673);
  not NOT_8476(g32882,g31376);
  not NOT_8477(g32883,g30735);
  not NOT_8478(g32884,g30825);
  not NOT_8479(g32885,g31021);
  not NOT_8480(g32886,g31327);
  not NOT_8481(g32887,g30614);
  not NOT_8482(g32888,g30673);
  not NOT_8483(g32889,g31376);
  not NOT_8484(g32890,g30735);
  not NOT_8485(g32891,g30825);
  not NOT_8486(g32892,g31021);
  not NOT_8487(g32893,g30937);
  not NOT_8488(g32894,g30614);
  not NOT_8489(g32895,g30673);
  not NOT_8490(g32896,g31376);
  not NOT_8491(g32897,g30735);
  not NOT_8492(g32898,g30825);
  not NOT_8493(g32899,g31021);
  not NOT_8494(g32900,g30937);
  not NOT_8495(g32901,g31327);
  not NOT_8496(g32902,g30673);
  not NOT_8497(g32903,g31376);
  not NOT_8498(g32904,g30735);
  not NOT_8499(g32905,g30825);
  not NOT_8500(g32906,g31021);
  not NOT_8501(g32907,g30937);
  not NOT_8502(g32908,g31327);
  not NOT_8503(g32909,g30614);
  not NOT_8504(g32911,g31376);
  not NOT_8505(g32912,g30735);
  not NOT_8506(g32913,g30825);
  not NOT_8507(g32914,g31672);
  not NOT_8508(g32915,g31710);
  not NOT_8509(g32916,g31021);
  not NOT_8510(g32917,g30937);
  not NOT_8511(g32918,g31327);
  not NOT_8512(g32919,g30735);
  not NOT_8513(g32920,g30825);
  not NOT_8514(g32921,g31672);
  not NOT_8515(g32922,g31710);
  not NOT_8516(g32923,g31021);
  not NOT_8517(g32924,g30937);
  not NOT_8518(g32925,g31327);
  not NOT_8519(g32926,g31376);
  not NOT_8520(g32927,g30825);
  not NOT_8521(g32928,g31672);
  not NOT_8522(g32929,g31710);
  not NOT_8523(g32930,g31021);
  not NOT_8524(g32931,g30937);
  not NOT_8525(g32932,g31327);
  not NOT_8526(g32933,g31376);
  not NOT_8527(g32934,g30735);
  not NOT_8528(g32935,g31672);
  not NOT_8529(g32936,g31710);
  not NOT_8530(g32937,g31021);
  not NOT_8531(g32938,g30937);
  not NOT_8532(g32939,g31327);
  not NOT_8533(g32940,g31376);
  not NOT_8534(g32941,g30735);
  not NOT_8535(g32942,g30825);
  not NOT_8536(g32943,g31710);
  not NOT_8537(g32944,g31021);
  not NOT_8538(g32945,g30937);
  not NOT_8539(g32946,g31327);
  not NOT_8540(g32947,g31376);
  not NOT_8541(g32948,g30735);
  not NOT_8542(g32949,g30825);
  not NOT_8543(g32950,g31672);
  not NOT_8544(g32951,g31021);
  not NOT_8545(g32952,g30937);
  not NOT_8546(g32953,g31327);
  not NOT_8547(g32954,g31376);
  not NOT_8548(g32955,g30735);
  not NOT_8549(g32956,g30825);
  not NOT_8550(g32957,g31672);
  not NOT_8551(g32958,g31710);
  not NOT_8552(g32959,g30937);
  not NOT_8553(g32960,g31327);
  not NOT_8554(g32961,g31376);
  not NOT_8555(g32962,g30735);
  not NOT_8556(g32963,g30825);
  not NOT_8557(g32964,g31672);
  not NOT_8558(g32965,g31710);
  not NOT_8559(g32966,g31021);
  not NOT_8560(g32967,g31327);
  not NOT_8561(g32968,g31376);
  not NOT_8562(g32969,g30735);
  not NOT_8563(g32970,g30825);
  not NOT_8564(g32971,g31672);
  not NOT_8565(g32972,g31710);
  not NOT_8566(g32973,g31021);
  not NOT_8567(g32974,g30937);
  not NOT_8568(I30537,g32027);
  not NOT_8569(g32975,I30537);
  not NOT_8570(g33072,g31945);
  not NOT_8571(I30641,g32024);
  not NOT_8572(g33079,I30641);
  not NOT_8573(I30644,g32024);
  not NOT_8574(g33080,I30644);
  not NOT_8575(I30686,g32381);
  not NOT_8576(g33120,I30686);
  not NOT_8577(g33127,g31950);
  not NOT_8578(g33136,g32057);
  not NOT_8579(g33142,g32072);
  not NOT_8580(I30766,g32363);
  not NOT_8581(g33228,I30766);
  not NOT_8582(g33246,g32212);
  not NOT_8583(g33250,g32186);
  not NOT_8584(g33258,g32296);
  not NOT_8585(g33326,g32318);
  not NOT_8586(I30861,g32383);
  not NOT_8587(g33335,I30861);
  not NOT_8588(g33346,g32132);
  not NOT_8589(g33354,g32329);
  not NOT_8590(g33375,g32377);
  not NOT_8591(I30901,g32407);
  not NOT_8592(g33377,I30901);
  not NOT_8593(I30904,g32424);
  not NOT_8594(g33378,I30904);
  not NOT_8595(g33382,g32033);
  not NOT_8596(g33385,g32038);
  not NOT_8597(g33388,g32382);
  not NOT_8598(g33391,g32384);
  not NOT_8599(g33413,g31971);
  not NOT_8600(g33424,g32415);
  not NOT_8601(g33426,g32017);
  not NOT_8602(g33430,g32421);
  not NOT_8603(I30959,g32021);
  not NOT_8604(g33435,I30959);
  not NOT_8605(I30962,g32021);
  not NOT_8606(g33436,I30962);
  not NOT_8607(g33442,g31937);
  not NOT_8608(I30971,g32015);
  not NOT_8609(g33443,I30971);
  not NOT_8610(g33451,g32132);
  not NOT_8611(I30980,g32132);
  not NOT_8612(g33454,I30980);
  not NOT_8613(I30983,g32433);
  not NOT_8614(g33455,I30983);
  not NOT_8615(I30986,g32437);
  not NOT_8616(g33456,I30986);
  not NOT_8617(I30989,g32441);
  not NOT_8618(g33457,I30989);
  not NOT_8619(I30992,g32445);
  not NOT_8620(g33458,I30992);
  not NOT_8621(I30995,g32449);
  not NOT_8622(g33459,I30995);
  not NOT_8623(I30998,g32453);
  not NOT_8624(g33460,I30998);
  not NOT_8625(I31361,g33120);
  not NOT_8626(g33533,I31361);
  not NOT_8627(I31459,g33219);
  not NOT_8628(g33631,I31459);
  not NOT_8629(g33635,g33436);
  not NOT_8630(I31463,g33318);
  not NOT_8631(g33636,I31463);
  not NOT_8632(I31466,g33318);
  not NOT_8633(g33637,I31466);
  not NOT_8634(I31469,g33388);
  not NOT_8635(g33638,I31469);
  not NOT_8636(I31474,g33212);
  not NOT_8637(g33641,I31474);
  not NOT_8638(I31477,g33391);
  not NOT_8639(g33645,I31477);
  not NOT_8640(I31482,g33204);
  not NOT_8641(g33648,I31482);
  not NOT_8642(I31486,g33197);
  not NOT_8643(g33653,I31486);
  not NOT_8644(g33658,g33080);
  not NOT_8645(I31491,g33283);
  not NOT_8646(g33659,I31491);
  not NOT_8647(I31494,g33283);
  not NOT_8648(g33660,I31494);
  not NOT_8649(I31497,g33187);
  not NOT_8650(g33661,I31497);
  not NOT_8651(I31500,g33176);
  not NOT_8652(g33665,I31500);
  not NOT_8653(I31504,g33164);
  not NOT_8654(g33670,I31504);
  not NOT_8655(I31515,g33187);
  not NOT_8656(g33682,I31515);
  not NOT_8657(g33686,g33187);
  not NOT_8658(I31523,g33187);
  not NOT_8659(g33688,I31523);
  not NOT_8660(I31528,g33219);
  not NOT_8661(g33691,I31528);
  not NOT_8662(g33695,g33187);
  not NOT_8663(I31535,g33377);
  not NOT_8664(g33696,I31535);
  not NOT_8665(I31539,g33212);
  not NOT_8666(g33698,I31539);
  not NOT_8667(I31545,g33219);
  not NOT_8668(g33702,I31545);
  not NOT_8669(I31550,g33204);
  not NOT_8670(g33705,I31550);
  not NOT_8671(I31555,g33212);
  not NOT_8672(g33708,I31555);
  not NOT_8673(I31561,g33197);
  not NOT_8674(g33712,I31561);
  not NOT_8675(I31564,g33204);
  not NOT_8676(g33713,I31564);
  not NOT_8677(I31569,g33197);
  not NOT_8678(g33716,I31569);
  not NOT_8679(I31581,g33164);
  not NOT_8680(g33726,I31581);
  not NOT_8681(I31586,g33149);
  not NOT_8682(g33729,I31586);
  not NOT_8683(I31597,g33187);
  not NOT_8684(g33736,I31597);
  not NOT_8685(I31604,g33176);
  not NOT_8686(g33744,I31604);
  not NOT_8687(I31607,g33164);
  not NOT_8688(g33750,I31607);
  not NOT_8689(I31610,g33149);
  not NOT_8690(g33755,I31610);
  not NOT_8691(I31616,g33219);
  not NOT_8692(g33761,I31616);
  not NOT_8693(I31619,g33212);
  not NOT_8694(g33766,I31619);
  not NOT_8695(I31622,g33204);
  not NOT_8696(g33772,I31622);
  not NOT_8697(I31625,g33197);
  not NOT_8698(g33778,I31625);
  not NOT_8699(g33797,g33306);
  not NOT_8700(g33799,g33299);
  not NOT_8701(I31642,g33204);
  not NOT_8702(g33800,I31642);
  not NOT_8703(g33804,g33250);
  not NOT_8704(I31650,g33212);
  not NOT_8705(g33806,I31650);
  not NOT_8706(I31659,g33219);
  not NOT_8707(g33813,I31659);
  not NOT_8708(I31672,g33149);
  not NOT_8709(g33827,I31672);
  not NOT_8710(I31686,g33164);
  not NOT_8711(g33839,I31686);
  not NOT_8712(I31694,g33176);
  not NOT_8713(g33845,I31694);
  not NOT_8714(I31701,g33164);
  not NOT_8715(g33850,I31701);
  not NOT_8716(I31724,g33076);
  not NOT_8717(g33874,I31724);
  not NOT_8718(I31727,g33076);
  not NOT_8719(g33875,I31727);
  not NOT_8720(g33888,g33346);
  not NOT_8721(I31748,g33228);
  not NOT_8722(g33894,I31748);
  not NOT_8723(I31751,g33228);
  not NOT_8724(g33895,I31751);
  not NOT_8725(I31770,g33197);
  not NOT_8726(g33912,I31770);
  not NOT_8727(I31776,g33204);
  not NOT_8728(g33916,I31776);
  not NOT_8729(I31779,g33212);
  not NOT_8730(g33917,I31779);
  not NOT_8731(I31782,g33219);
  not NOT_8732(g33918,I31782);
  not NOT_8733(I31786,g33197);
  not NOT_8734(g33920,I31786);
  not NOT_8735(I31791,g33354);
  not NOT_8736(g33923,I31791);
  not NOT_8737(I31796,g33176);
  not NOT_8738(g33926,I31796);
  not NOT_8739(I31800,g33164);
  not NOT_8740(g33928,I31800);
  not NOT_8741(I31803,g33176);
  not NOT_8742(g33929,I31803);
  not NOT_8743(I31807,g33149);
  not NOT_8744(g33931,I31807);
  not NOT_8745(I31810,g33164);
  not NOT_8746(g33932,I31810);
  not NOT_8747(I31814,g33149);
  not NOT_8748(g33934,I31814);
  not NOT_8749(I31817,g33323);
  not NOT_8750(g33935,I31817);
  not NOT_8751(I31820,g33323);
  not NOT_8752(g33936,I31820);
  not NOT_8753(I31823,g33149);
  not NOT_8754(g33937,I31823);
  not NOT_8755(I31829,g33454);
  not NOT_8756(g33944,I31829);
  not NOT_8757(I31878,g33696);
  not NOT_8758(g33959,I31878);
  not NOT_8759(g34042,g33674);
  not NOT_8760(g34044,g33675);
  not NOT_8761(g34047,g33637);
  not NOT_8762(g34049,g33678);
  not NOT_8763(g34052,g33635);
  not NOT_8764(g34053,g33683);
  not NOT_8765(g34058,g33660);
  not NOT_8766(g34059,g33658);
  not NOT_8767(g34060,g33704);
  not NOT_8768(g34062,g33711);
  not NOT_8769(g34068,g33728);
  not NOT_8770(g34070,g33725);
  not NOT_8771(g34094,g33772);
  not NOT_8772(I32051,g33631);
  not NOT_8773(g34118,I32051);
  not NOT_8774(I32056,g33641);
  not NOT_8775(g34121,I32056);
  not NOT_8776(I32059,g33648);
  not NOT_8777(g34122,I32059);
  not NOT_8778(I32062,g33653);
  not NOT_8779(g34123,I32062);
  not NOT_8780(g34124,g33819);
  not NOT_8781(I32067,g33661);
  not NOT_8782(g34126,I32067);
  not NOT_8783(I32071,g33665);
  not NOT_8784(g34130,I32071);
  not NOT_8785(I32074,g33670);
  not NOT_8786(g34131,I32074);
  not NOT_8787(g34132,g33831);
  not NOT_8788(I32079,g33937);
  not NOT_8789(g34134,I32079);
  not NOT_8790(I32089,g33665);
  not NOT_8791(g34142,I32089);
  not NOT_8792(I32093,g33670);
  not NOT_8793(g34144,I32093);
  not NOT_8794(I32096,g33641);
  not NOT_8795(g34145,I32096);
  not NOT_8796(g34147,g33823);
  not NOT_8797(I32103,g33661);
  not NOT_8798(g34150,I32103);
  not NOT_8799(I32106,g33653);
  not NOT_8800(g34151,I32106);
  not NOT_8801(I32109,g33631);
  not NOT_8802(g34152,I32109);
  not NOT_8803(g34156,g33907);
  not NOT_8804(I32116,g33937);
  not NOT_8805(g34159,I32116);
  not NOT_8806(I32119,g33648);
  not NOT_8807(g34160,I32119);
  not NOT_8808(g34161,g33851);
  not NOT_8809(g34181,g33913);
  not NOT_8810(g34188,g33875);
  not NOT_8811(g34192,g33921);
  not NOT_8812(I32150,g33923);
  not NOT_8813(g34195,I32150);
  not NOT_8814(g34197,g33812);
  not NOT_8815(g34200,g33895);
  not NOT_8816(I32158,g33791);
  not NOT_8817(g34201,I32158);
  not NOT_8818(I32161,g33791);
  not NOT_8819(g34202,I32161);
  not NOT_8820(g34208,g33838);
  not NOT_8821(I32170,g33638);
  not NOT_8822(g34209,I32170);
  not NOT_8823(I32173,g33645);
  not NOT_8824(g34210,I32173);
  not NOT_8825(I32192,g33628);
  not NOT_8826(g34221,I32192);
  not NOT_8827(I32195,g33628);
  not NOT_8828(g34222,I32195);
  not NOT_8829(g34229,g33936);
  not NOT_8830(I32222,g34118);
  not NOT_8831(g34241,I32222);
  not NOT_8832(I32225,g34121);
  not NOT_8833(g34242,I32225);
  not NOT_8834(I32228,g34122);
  not NOT_8835(g34243,I32228);
  not NOT_8836(I32231,g34123);
  not NOT_8837(g34244,I32231);
  not NOT_8838(I32234,g34126);
  not NOT_8839(g34245,I32234);
  not NOT_8840(I32237,g34130);
  not NOT_8841(g34246,I32237);
  not NOT_8842(I32240,g34131);
  not NOT_8843(g34247,I32240);
  not NOT_8844(I32243,g34134);
  not NOT_8845(g34248,I32243);
  not NOT_8846(g34270,g34159);
  not NOT_8847(g34271,g34160);
  not NOT_8848(g34272,g34229);
  not NOT_8849(g34275,g34047);
  not NOT_8850(g34276,g34058);
  not NOT_8851(I32274,g34195);
  not NOT_8852(g34277,I32274);
  not NOT_8853(I32284,g34052);
  not NOT_8854(g34285,I32284);
  not NOT_8855(I32297,g34059);
  not NOT_8856(g34296,I32297);
  not NOT_8857(g34299,g34080);
  not NOT_8858(I32305,g34209);
  not NOT_8859(g34302,I32305);
  not NOT_8860(I32309,g34210);
  not NOT_8861(g34304,I32309);
  not NOT_8862(g34307,g34087);
  not NOT_8863(g34308,g34088);
  not NOT_8864(g34311,g34097);
  not NOT_8865(g34312,g34098);
  not NOT_8866(g34313,g34086);
  not NOT_8867(g34315,g34085);
  not NOT_8868(g34316,g34093);
  not NOT_8869(g34317,g34115);
  not NOT_8870(g34320,g34119);
  not NOT_8871(g34323,g34105);
  not NOT_8872(g34325,g34092);
  not NOT_8873(g34326,g34091);
  not NOT_8874(g34327,g34108);
  not NOT_8875(g34328,g34096);
  not NOT_8876(g34336,g34112);
  not NOT_8877(g34339,g34077);
  not NOT_8878(g34343,g34089);
  not NOT_8879(I32352,g34169);
  not NOT_8880(g34345,I32352);
  not NOT_8881(g34346,g34162);
  not NOT_8882(g34351,g34174);
  not NOT_8883(I32364,g34208);
  not NOT_8884(g34358,I32364);
  not NOT_8885(I32388,g34153);
  not NOT_8886(g34383,I32388);
  not NOT_8887(I32391,g34153);
  not NOT_8888(g34384,I32391);
  not NOT_8889(g34387,g34188);
  not NOT_8890(g34391,g34200);
  not NOT_8891(g34392,g34202);
  not NOT_8892(g34400,g34142);
  not NOT_8893(g34408,g34144);
  not NOT_8894(g34409,g34145);
  not NOT_8895(g34418,g34150);
  not NOT_8896(g34419,g34151);
  not NOT_8897(g34420,g34152);
  not NOT_8898(g34423,g34222);
  not NOT_8899(I32446,g34127);
  not NOT_8900(g34425,I32446);
  not NOT_8901(I32449,g34127);
  not NOT_8902(g34426,I32449);
  not NOT_8903(I32452,g34241);
  not NOT_8904(g34427,I32452);
  not NOT_8905(I32455,g34242);
  not NOT_8906(g34428,I32455);
  not NOT_8907(I32458,g34243);
  not NOT_8908(g34429,I32458);
  not NOT_8909(I32461,g34244);
  not NOT_8910(g34430,I32461);
  not NOT_8911(I32464,g34245);
  not NOT_8912(g34431,I32464);
  not NOT_8913(I32467,g34246);
  not NOT_8914(g34432,I32467);
  not NOT_8915(I32470,g34247);
  not NOT_8916(g34433,I32470);
  not NOT_8917(I32473,g34248);
  not NOT_8918(g34434,I32473);
  not NOT_8919(I32476,g34277);
  not NOT_8920(g34435,I32476);
  not NOT_8921(I32479,g34302);
  not NOT_8922(g34436,I32479);
  not NOT_8923(I32482,g34304);
  not NOT_8924(g34437,I32482);
  not NOT_8925(g34471,g34423);
  not NOT_8926(I32525,g34285);
  not NOT_8927(g34472,I32525);
  not NOT_8928(g34473,g34426);
  not NOT_8929(I32535,g34296);
  not NOT_8930(g34480,I32535);
  not NOT_8931(I32547,g34397);
  not NOT_8932(g34490,I32547);
  not NOT_8933(I32550,g34398);
  not NOT_8934(g34491,I32550);
  not NOT_8935(g34501,g34400);
  not NOT_8936(g34504,g34408);
  not NOT_8937(g34505,g34409);
  not NOT_8938(g34510,g34418);
  not NOT_8939(g34511,g34419);
  not NOT_8940(g34512,g34420);
  not NOT_8941(g34521,g34270);
  not NOT_8942(g34522,g34271);
  not NOT_8943(I32591,g34287);
  not NOT_8944(g34530,I32591);
  not NOT_8945(I32594,g34298);
  not NOT_8946(g34531,I32594);
  not NOT_8947(I32601,g34319);
  not NOT_8948(g34536,I32601);
  not NOT_8949(g34539,g34354);
  not NOT_8950(I32607,g34358);
  not NOT_8951(g34540,I32607);
  not NOT_8952(g34543,g34359);
  not NOT_8953(I32613,g34329);
  not NOT_8954(g34544,I32613);
  not NOT_8955(I32617,g34333);
  not NOT_8956(g34549,I32617);
  not NOT_8957(I32621,g34335);
  not NOT_8958(g34553,I32621);
  not NOT_8959(g34559,g34384);
  not NOT_8960(I32639,g34345);
  not NOT_8961(g34569,I32639);
  not NOT_8962(g34570,g34392);
  not NOT_8963(I32645,g34367);
  not NOT_8964(g34573,I32645);
  not NOT_8965(I32648,g34371);
  not NOT_8966(g34574,I32648);
  not NOT_8967(I32651,g34375);
  not NOT_8968(g34575,I32651);
  not NOT_8969(I32654,g34378);
  not NOT_8970(g34576,I32654);
  not NOT_8971(I32659,g34391);
  not NOT_8972(g34579,I32659);
  not NOT_8973(I32665,g34386);
  not NOT_8974(g34583,I32665);
  not NOT_8975(I32671,g34388);
  not NOT_8976(g34587,I32671);
  not NOT_8977(I32675,g34427);
  not NOT_8978(g34589,I32675);
  not NOT_8979(I32678,g34428);
  not NOT_8980(g34590,I32678);
  not NOT_8981(I32681,g34429);
  not NOT_8982(g34591,I32681);
  not NOT_8983(I32684,g34430);
  not NOT_8984(g34592,I32684);
  not NOT_8985(I32687,g34431);
  not NOT_8986(g34593,I32687);
  not NOT_8987(I32690,g34432);
  not NOT_8988(g34594,I32690);
  not NOT_8989(I32693,g34433);
  not NOT_8990(g34595,I32693);
  not NOT_8991(I32696,g34434);
  not NOT_8992(g34596,I32696);
  not NOT_8993(I32699,g34569);
  not NOT_8994(g34597,I32699);
  not NOT_8995(I32752,g34510);
  not NOT_8996(g34648,I32752);
  not NOT_8997(I32763,g34511);
  not NOT_8998(g34653,I32763);
  not NOT_8999(I32766,g34522);
  not NOT_9000(g34654,I32766);
  not NOT_9001(I32770,g34505);
  not NOT_9002(g34656,I32770);
  not NOT_9003(I32775,g34512);
  not NOT_9004(g34659,I32775);
  not NOT_9005(g34660,g34473);
  not NOT_9006(I32782,g34571);
  not NOT_9007(g34664,I32782);
  not NOT_9008(I32788,g34577);
  not NOT_9009(g34668,I32788);
  not NOT_9010(I32791,g34578);
  not NOT_9011(g34669,I32791);
  not NOT_9012(I32794,g34580);
  not NOT_9013(g34670,I32794);
  not NOT_9014(I32797,g34581);
  not NOT_9015(g34671,I32797);
  not NOT_9016(I32800,g34582);
  not NOT_9017(g34672,I32800);
  not NOT_9018(I32803,g34584);
  not NOT_9019(g34673,I32803);
  not NOT_9020(I32806,g34585);
  not NOT_9021(g34674,I32806);
  not NOT_9022(I32809,g34586);
  not NOT_9023(g34675,I32809);
  not NOT_9024(I32812,g34588);
  not NOT_9025(g34676,I32812);
  not NOT_9026(I32815,g34470);
  not NOT_9027(g34677,I32815);
  not NOT_9028(I32820,g34474);
  not NOT_9029(g34680,I32820);
  not NOT_9030(I32824,g34475);
  not NOT_9031(g34682,I32824);
  not NOT_9032(I32827,g34477);
  not NOT_9033(g34683,I32827);
  not NOT_9034(I32834,g34472);
  not NOT_9035(g34688,I32834);
  not NOT_9036(I32837,g34498);
  not NOT_9037(g34689,I32837);
  not NOT_9038(I32840,g34480);
  not NOT_9039(g34690,I32840);
  not NOT_9040(I32843,g34499);
  not NOT_9041(g34691,I32843);
  not NOT_9042(I32846,g34502);
  not NOT_9043(g34692,I32846);
  not NOT_9044(g34697,g34545);
  not NOT_9045(g34698,g34550);
  not NOT_9046(I32855,g34540);
  not NOT_9047(g34699,I32855);
  not NOT_9048(g34711,g34559);
  not NOT_9049(I32868,g34579);
  not NOT_9050(g34712,I32868);
  not NOT_9051(I32871,g34521);
  not NOT_9052(g34713,I32871);
  not NOT_9053(I32874,g34504);
  not NOT_9054(g34714,I32874);
  not NOT_9055(I32878,g34501);
  not NOT_9056(g34716,I32878);
  not NOT_9057(I32881,g34688);
  not NOT_9058(g34717,I32881);
  not NOT_9059(I32884,g34690);
  not NOT_9060(g34718,I32884);
  not NOT_9061(I32904,g34708);
  not NOT_9062(g34736,I32904);
  not NOT_9063(I32909,g34712);
  not NOT_9064(g34739,I32909);
  not NOT_9065(I32921,g34650);
  not NOT_9066(g34749,I32921);
  not NOT_9067(I32929,g34649);
  not NOT_9068(g34755,I32929);
  not NOT_9069(I32935,g34657);
  not NOT_9070(g34759,I32935);
  not NOT_9071(I32938,g34663);
  not NOT_9072(g34760,I32938);
  not NOT_9073(g34766,g34703);
  not NOT_9074(I32947,g34659);
  not NOT_9075(g34767,I32947);
  not NOT_9076(I32950,g34713);
  not NOT_9077(g34768,I32950);
  not NOT_9078(I32953,g34656);
  not NOT_9079(g34769,I32953);
  not NOT_9080(I32956,g34654);
  not NOT_9081(g34770,I32956);
  not NOT_9082(I32960,g34653);
  not NOT_9083(g34772,I32960);
  not NOT_9084(I32963,g34650);
  not NOT_9085(g34773,I32963);
  not NOT_9086(I32967,g34648);
  not NOT_9087(g34775,I32967);
  not NOT_9088(I32970,g34716);
  not NOT_9089(g34776,I32970);
  not NOT_9090(I32973,g34714);
  not NOT_9091(g34777,I32973);
  not NOT_9092(I32976,g34699);
  not NOT_9093(g34778,I32976);
  not NOT_9094(I32982,g34749);
  not NOT_9095(g34784,I32982);
  not NOT_9096(I32985,g34736);
  not NOT_9097(g34785,I32985);
  not NOT_9098(I32988,g34755);
  not NOT_9099(g34786,I32988);
  not NOT_9100(I32991,g34759);
  not NOT_9101(g34787,I32991);
  not NOT_9102(I32994,g34739);
  not NOT_9103(g34788,I32994);
  not NOT_9104(I32997,g34760);
  not NOT_9105(g34789,I32997);
  not NOT_9106(I33020,g34781);
  not NOT_9107(g34810,I33020);
  not NOT_9108(I33024,g34783);
  not NOT_9109(g34812,I33024);
  not NOT_9110(I33027,g34767);
  not NOT_9111(g34813,I33027);
  not NOT_9112(I33030,g34768);
  not NOT_9113(g34816,I33030);
  not NOT_9114(I33034,g34769);
  not NOT_9115(g34820,I33034);
  not NOT_9116(I33037,g34770);
  not NOT_9117(g34823,I33037);
  not NOT_9118(I33041,g34772);
  not NOT_9119(g34827,I33041);
  not NOT_9120(I33044,g34775);
  not NOT_9121(g34830,I33044);
  not NOT_9122(I33047,g34776);
  not NOT_9123(g34833,I33047);
  not NOT_9124(I33050,g34777);
  not NOT_9125(g34836,I33050);
  not NOT_9126(I33053,g34778);
  not NOT_9127(g34839,I33053);
  not NOT_9128(I33056,g34778);
  not NOT_9129(g34840,I33056);
  not NOT_9130(g34844,g34737);
  not NOT_9131(g34845,g34773);
  not NOT_9132(I33064,g34784);
  not NOT_9133(g34846,I33064);
  not NOT_9134(I33067,g34812);
  not NOT_9135(g34847,I33067);
  not NOT_9136(I33070,g34810);
  not NOT_9137(g34848,I33070);
  not NOT_9138(I33075,g34843);
  not NOT_9139(g34851,I33075);
  not NOT_9140(g34852,g34845);
  not NOT_9141(I33079,g34809);
  not NOT_9142(g34855,I33079);
  not NOT_9143(g34864,g34840);
  not NOT_9144(I33103,g34846);
  not NOT_9145(g34877,I33103);
  not NOT_9146(I33106,g34855);
  not NOT_9147(g34878,I33106);
  not NOT_9148(I33109,g34851);
  not NOT_9149(g34879,I33109);
  not NOT_9150(g34883,g34852);
  not NOT_9151(I33119,g34852);
  not NOT_9152(g34893,I33119);
  not NOT_9153(g34910,g34864);
  not NOT_9154(I33131,g34906);
  not NOT_9155(g34913,I33131);
  not NOT_9156(I33134,g34906);
  not NOT_9157(g34914,I33134);
  not NOT_9158(I33137,g34884);
  not NOT_9159(g34915,I33137);
  not NOT_9160(I33140,g34884);
  not NOT_9161(g34916,I33140);
  not NOT_9162(I33143,g34903);
  not NOT_9163(g34917,I33143);
  not NOT_9164(I33146,g34903);
  not NOT_9165(g34918,I33146);
  not NOT_9166(I33149,g34900);
  not NOT_9167(g34919,I33149);
  not NOT_9168(I33152,g34900);
  not NOT_9169(g34920,I33152);
  not NOT_9170(I33155,g34897);
  not NOT_9171(g34921,I33155);
  not NOT_9172(I33158,g34897);
  not NOT_9173(g34922,I33158);
  not NOT_9174(I33161,g34894);
  not NOT_9175(g34923,I33161);
  not NOT_9176(I33164,g34894);
  not NOT_9177(g34924,I33164);
  not NOT_9178(I33167,g34890);
  not NOT_9179(g34925,I33167);
  not NOT_9180(I33170,g34890);
  not NOT_9181(g34926,I33170);
  not NOT_9182(I33173,g34887);
  not NOT_9183(g34927,I33173);
  not NOT_9184(I33176,g34887);
  not NOT_9185(g34928,I33176);
  not NOT_9186(I33179,g34893);
  not NOT_9187(g34929,I33179);
  not NOT_9188(I33182,g34910);
  not NOT_9189(g34930,I33182);
  not NOT_9190(g34932,g34914);
  not NOT_9191(g34933,g34916);
  not NOT_9192(g34934,g34918);
  not NOT_9193(I33189,g34929);
  not NOT_9194(g34935,I33189);
  not NOT_9195(g34938,g34920);
  not NOT_9196(g34939,g34922);
  not NOT_9197(g34940,g34924);
  not NOT_9198(g34941,g34926);
  not NOT_9199(g34942,g34928);
  not NOT_9200(I33197,g34930);
  not NOT_9201(g34943,I33197);
  not NOT_9202(g34944,g34932);
  not NOT_9203(g34945,g34933);
  not NOT_9204(g34946,g34934);
  not NOT_9205(g34947,g34938);
  not NOT_9206(g34949,g34939);
  not NOT_9207(g34950,g34940);
  not NOT_9208(g34951,g34941);
  not NOT_9209(g34952,g34942);
  not NOT_9210(I33210,g34943);
  not NOT_9211(g34954,I33210);
  not NOT_9212(I33214,g34954);
  not NOT_9213(g34956,I33214);
  not NOT_9214(I33218,g34955);
  not NOT_9215(g34960,I33218);
  not NOT_9216(I33232,g34957);
  not NOT_9217(g34972,I33232);
  not NOT_9218(I33235,g34957);
  not NOT_9219(g34973,I33235);
  not NOT_9220(g34981,g34973);
  not NOT_9221(I33246,g34970);
  not NOT_9222(g34982,I33246);
  not NOT_9223(I33249,g34971);
  not NOT_9224(g34983,I33249);
  not NOT_9225(I33252,g34974);
  not NOT_9226(g34984,I33252);
  not NOT_9227(I33255,g34975);
  not NOT_9228(g34985,I33255);
  not NOT_9229(I33258,g34976);
  not NOT_9230(g34986,I33258);
  not NOT_9231(I33261,g34977);
  not NOT_9232(g34987,I33261);
  not NOT_9233(I33264,g34978);
  not NOT_9234(g34988,I33264);
  not NOT_9235(I33267,g34979);
  not NOT_9236(g34989,I33267);
  not NOT_9237(I33270,g34982);
  not NOT_9238(g34990,I33270);
  not NOT_9239(I33273,g34984);
  not NOT_9240(g34991,I33273);
  not NOT_9241(I33276,g34985);
  not NOT_9242(g34992,I33276);
  not NOT_9243(I33279,g34986);
  not NOT_9244(g34993,I33279);
  not NOT_9245(I33282,g34987);
  not NOT_9246(g34994,I33282);
  not NOT_9247(I33285,g34988);
  not NOT_9248(g34995,I33285);
  not NOT_9249(I33288,g34989);
  not NOT_9250(g34996,I33288);
  not NOT_9251(I33291,g34983);
  not NOT_9252(g34997,I33291);
  not NOT_9253(g34998,g34981);
  not NOT_9254(I33297,g35000);
  not NOT_9255(g35001,I33297);
  not NOT_9256(I33300,g35001);
  not NOT_9257(g35002,I33300);
  and AND_9258(g7251,g452,g392);
  and AND_9259(g7396,g392,g441);
  and AND_9260(g7469,g4382,g4438);
  and AND_9261(g7511,g2145,g2138,g2130);
  and AND_9262(g7520,g2704,g2697,g2689);
  and AND_9263(g7685,g4382,g4375);
  and AND_9264(g7696,g2955,g2950);
  and AND_9265(g7763,g2965,g2960);
  and AND_9266(g7777,g723,g822,g817);
  and AND_9267(g7804,g2975,g2970);
  and AND_9268(g7918,g1205,g1087);
  and AND_9269(g7948,g1548,g1430);
  and AND_9270(g8234,g4515,g4521);
  and AND_9271(g8530,g2902,g2907);
  and AND_9272(g8583,g2917,g2912);
  and AND_9273(g8643,g2927,g2922);
  and AND_9274(g8690,g2941,g2936);
  and AND_9275(g8721,g385,g376,g365);
  and AND_9276(g9217,g632,g626);
  and AND_9277(g9479,g305,g324);
  and AND_9278(g9906,g996,g1157);
  and AND_9279(g9967,g1178,g1157);
  and AND_9280(g9968,g1339,g1500);
  and AND_9281(g10034,g1521,g1500);
  and AND_9282(g10290,g4358,g4349);
  and AND_9283(I13862,g7232,g7219,g7258);
  and AND_9284(g10476,g7244,g7259,I13862);
  and AND_9285(g10501,g1233,g9007);
  and AND_9286(g10528,g1576,g9051);
  and AND_9287(g10543,g8238,g437);
  and AND_9288(g10565,g8182,g424);
  and AND_9289(g10588,g7004,g5297);
  and AND_9290(I13937,g7340,g7293,g7261);
  and AND_9291(g10590,g7246,g7392,I13937);
  and AND_9292(g10616,g7998,g174);
  and AND_9293(g10619,g3080,g7907);
  and AND_9294(g10624,g8387,g3072);
  and AND_9295(g10625,g3431,g7926);
  and AND_9296(g10626,g4057,g7927);
  and AND_9297(g10632,g7475,g7441,g890);
  and AND_9298(g10654,g3085,g8434);
  and AND_9299(g10655,g8440,g3423);
  and AND_9300(g10656,g3782,g7952);
  and AND_9301(g10657,g8451,g4064);
  and AND_9302(g10665,g209,g8292);
  and AND_9303(g10674,g6841,g10200,g2130);
  and AND_9304(g10675,g3436,g8500);
  and AND_9305(g10676,g8506,g3774);
  and AND_9306(g10677,g4141,g7611);
  and AND_9307(g10683,g7289,g4438);
  and AND_9308(g10684,g7998,g411);
  and AND_9309(g10704,g2145,g10200,g2130);
  and AND_9310(g10705,g6850,g10219,g2689);
  and AND_9311(g10706,g3338,g8691);
  and AND_9312(g10707,g3787,g8561);
  and AND_9313(g10719,g6841,g2138,g2130);
  and AND_9314(g10720,g2704,g10219,g2689);
  and AND_9315(g10721,g3288,g6875,g3274,g8481);
  and AND_9316(g10724,g3689,g8728);
  and AND_9317(g10732,g6850,g2697,g2689);
  and AND_9318(g10733,g3639,g6905,g3625,g8542);
  and AND_9319(g10736,g4040,g8751);
  and AND_9320(g10756,g3990,g6928,g3976,g8595);
  and AND_9321(g10822,g4264,g8514);
  and AND_9322(g10823,g7704,g5180,g5188);
  and AND_9323(g10827,g8914,g4258);
  and AND_9324(g10828,g6888,g7640);
  and AND_9325(g10829,g7289,g4375);
  and AND_9326(g10838,g7738,g5527,g5535);
  and AND_9327(g10841,g8509,g8567);
  and AND_9328(g10856,g4269,g8967);
  and AND_9329(g10869,g7766,g5873,g5881);
  and AND_9330(g10873,g3004,g9015);
  and AND_9331(g10874,g7791,g6219,g6227);
  and AND_9332(g10878,g7858,g1135);
  and AND_9333(g10883,g3355,g9061);
  and AND_9334(g10887,g7812,g6565,g6573);
  and AND_9335(g10890,g7858,g1105);
  and AND_9336(g10896,g1205,g8654);
  and AND_9337(g10898,g3706,g9100);
  and AND_9338(g10902,g7858,g1129);
  and AND_9339(g10917,g9174,g1087);
  and AND_9340(g10921,g1548,g8685);
  and AND_9341(g10925,g7858,g956);
  and AND_9342(g10934,g9197,g7918);
  and AND_9343(g10947,g9200,g1430);
  and AND_9344(g10948,g7880,g1478);
  and AND_9345(g10966,g9226,g7948);
  and AND_9346(g10967,g7880,g1448);
  and AND_9347(g10970,g854,g9582);
  and AND_9348(g10998,g8567,g8509,g8451,g7650);
  and AND_9349(g10999,g7880,g1472);
  and AND_9350(g11003,g7880,g1300);
  and AND_9351(g11010,g4698,g8933);
  and AND_9352(g11016,g4888,g8984);
  and AND_9353(g11018,g7655,g7643,g7627);
  and AND_9354(g11019,g5092,g9036);
  and AND_9355(g11023,g9669,g5084);
  and AND_9356(g11024,g5436,g9070);
  and AND_9357(g11027,g5097,g9724);
  and AND_9358(g11028,g9730,g5428);
  and AND_9359(g11029,g5782,g9103);
  and AND_9360(g11032,g9354,g7717);
  and AND_9361(g11035,g5441,g9800);
  and AND_9362(g11036,g9806,g5774);
  and AND_9363(g11037,g6128,g9184);
  and AND_9364(g11044,g5343,g10124);
  and AND_9365(g11045,g5787,g9883);
  and AND_9366(g11046,g9889,g6120);
  and AND_9367(g11047,g6474,g9212);
  and AND_9368(g11083,g8836,g802);
  and AND_9369(g11111,g5297,g7004,g5283,g9780);
  and AND_9370(g11114,g5689,g10160);
  and AND_9371(g11115,g6133,g9954);
  and AND_9372(g11116,g9960,g6466);
  and AND_9373(g11123,g5644,g7028,g5630,g9864);
  and AND_9374(g11126,g6035,g10185);
  and AND_9375(g11127,g6479,g10022);
  and AND_9376(g11139,g5990,g7051,g5976,g9935);
  and AND_9377(g11142,g6381,g10207);
  and AND_9378(I14198,g225,g8237,g232,g8180);
  and AND_9379(g11144,g239,g8136,g246,I14198);
  and AND_9380(g11160,g6336,g7074,g6322,g10003);
  and AND_9381(g11163,g6727,g10224);
  and AND_9382(I14225,g8457,g255,g8406,g262);
  and AND_9383(g11166,g8363,g269,g8296,I14225);
  and AND_9384(g11178,g6682,g7097,g6668,g10061);
  and AND_9385(g11205,g8217,g8439);
  and AND_9386(g11223,g8281,g8505);
  and AND_9387(g11244,g8346,g8566);
  and AND_9388(g11366,g5016,g10338);
  and AND_9389(g11397,g5360,g7139);
  and AND_9390(g11427,g5706,g7158);
  and AND_9391(g11449,g6052,g7175);
  and AND_9392(g11496,g4382,g7495);
  and AND_9393(g11497,g6398,g7192);
  and AND_9394(g11546,g7289,g4375);
  and AND_9395(g11740,g8769,g703);
  and AND_9396(g11890,g7499,g9155);
  and AND_9397(g11893,g1668,g7268);
  and AND_9398(g11915,g1802,g7315);
  and AND_9399(g11916,g2227,g7328);
  and AND_9400(g11937,g1936,g7362);
  and AND_9401(g11939,g2361,g7380);
  and AND_9402(g11956,g2070,g7411);
  and AND_9403(g11960,g2495,g7424);
  and AND_9404(g11967,g311,g7802);
  and AND_9405(g11978,g2629,g7462);
  and AND_9406(g12015,g1002,g7567);
  and AND_9407(g12027,g9499,g9729);
  and AND_9408(g12043,g1345,g7601);
  and AND_9409(g12065,g9557,g9805);
  and AND_9410(g12099,g9619,g9888);
  and AND_9411(g12135,g9684,g9959);
  and AND_9412(g12179,g9745,g10027);
  and AND_9413(g12186,g1178,g7519);
  and AND_9414(g12219,g1189,g7532);
  and AND_9415(g12220,g1521,g7535);
  and AND_9416(g12259,g9480,g640);
  and AND_9417(g12284,g1532,g7557);
  and AND_9418(g12527,g8680,g667);
  and AND_9419(g12641,g10295,g3171,g3179);
  and AND_9420(g12687,g9024,g8977);
  and AND_9421(g12692,g10323,g3522,g3530);
  and AND_9422(g12730,g9024,g4349);
  and AND_9423(g12735,g7121,g3873,g3881);
  and AND_9424(g12761,g969,g7567);
  and AND_9425(g12762,g4358,g8977);
  and AND_9426(g12794,g1008,g7567);
  and AND_9427(g12795,g1312,g7601);
  and AND_9428(g12812,g518,g9158);
  and AND_9429(g12817,g1351,g7601);
  and AND_9430(g12920,g1227,g10960);
  and AND_9431(g12924,g1570,g10980);
  and AND_9432(g12931,g392,g11048);
  and AND_9433(g12939,g405,g11048);
  and AND_9434(g12953,g411,g11048);
  and AND_9435(g12979,g424,g11048);
  and AND_9436(g13019,g194,g11737);
  and AND_9437(g13020,g401,g11048);
  and AND_9438(g13025,g8431,g11026);
  and AND_9439(g13029,g8359,g11030);
  and AND_9440(g13030,g429,g11048);
  and AND_9441(g13035,g8497,g11033);
  and AND_9442(g13038,g8509,g11034);
  and AND_9443(g13042,g433,g11048);
  and AND_9444(g13046,g6870,g11270);
  and AND_9445(g13047,g8534,g11042);
  and AND_9446(g13048,g8558,g11043);
  and AND_9447(g13059,g6900,g11303);
  and AND_9448(g13060,g8587,g11110);
  and AND_9449(g13063,g8567,g10808);
  and AND_9450(g13080,g6923,g11357);
  and AND_9451(g13081,g8626,g11122);
  and AND_9452(g13156,g10816,g10812,g10805);
  and AND_9453(g13221,g6946,g11425);
  and AND_9454(g13247,g8964,g11316);
  and AND_9455(g13252,g11561,g11511,g11469,g699);
  and AND_9456(g13265,g9018,g11493);
  and AND_9457(g13277,g3195,g11432);
  and AND_9458(g13282,g3546,g11480);
  and AND_9459(g13287,g1221,g11472);
  and AND_9460(g13290,g3897,g11534);
  and AND_9461(g13294,g1564,g11513);
  and AND_9462(g13299,g437,g11048);
  and AND_9463(g13306,g441,g11048);
  and AND_9464(g13313,g475,g11048);
  and AND_9465(g13319,g4076,g8812,g10658,g8757);
  and AND_9466(g13320,g417,g11048);
  and AND_9467(g13321,g847,g11048);
  and AND_9468(g13324,g854,g11326);
  and AND_9469(g13333,g4743,g11755);
  and AND_9470(g13345,g4754,g11773);
  and AND_9471(g13349,g4933,g11780);
  and AND_9472(g13383,g4765,g11797);
  and AND_9473(g13384,g4944,g11804);
  and AND_9474(g13393,g703,g11048);
  and AND_9475(g13411,g4955,g11834);
  and AND_9476(g13415,g837,g11048);
  and AND_9477(g13436,g9721,g11811);
  and AND_9478(g13461,g2719,g11819);
  and AND_9479(g13473,g9797,g11841);
  and AND_9480(g13491,g6999,g12160);
  and AND_9481(g13492,g9856,g11865);
  and AND_9482(g13493,g9880,g11866);
  and AND_9483(g13497,g2724,g12155);
  and AND_9484(g13507,g7023,g12198);
  and AND_9485(g13508,g9927,g11888);
  and AND_9486(g13509,g9951,g11889);
  and AND_9487(g13523,g7046,g12246);
  and AND_9488(g13524,g9995,g11910);
  and AND_9489(g13525,g10019,g11911);
  and AND_9490(g13541,g7069,g12308);
  and AND_9491(g13542,g10053,g11927);
  and AND_9492(g13564,g4480,g12820);
  and AND_9493(g13566,g7092,g12358);
  and AND_9494(g13567,g10102,g11948);
  and AND_9495(g13604,g4495,g10487);
  and AND_9496(g13632,g10232,g12228);
  and AND_9497(g13633,g4567,g10509);
  and AND_9498(g13656,g278,g11144);
  and AND_9499(g13671,g4498,g10532);
  and AND_9500(g13697,g11166,g8608);
  and AND_9501(g13737,g4501,g10571);
  and AND_9502(g13738,g8880,g10572);
  and AND_9503(I16111,g8691,g11409,g11381);
  and AND_9504(g13771,g11441,g11355,g11302,I16111);
  and AND_9505(g13778,g4540,g10597);
  and AND_9506(I16129,g8728,g11443,g11411);
  and AND_9507(g13805,g11489,g11394,g11356,I16129);
  and AND_9508(g13807,g4504,g10606);
  and AND_9509(g13808,g4543,g10607);
  and AND_9510(I16143,g8751,g11491,g11445);
  and AND_9511(g13830,g11543,g11424,g11395,I16143);
  and AND_9512(g13832,g8880,g10612);
  and AND_9513(g13833,g4546,g10613);
  and AND_9514(g13853,g4549,g10620);
  and AND_9515(g13887,g5204,g12402);
  and AND_9516(g13912,g5551,g12450);
  and AND_9517(g13942,g5897,g12512);
  and AND_9518(g13974,g6243,g12578);
  and AND_9519(g13998,g6589,g12629);
  and AND_9520(g14028,g8673,g11797);
  and AND_9521(g14035,g699,g11048);
  and AND_9522(g14061,g8715,g11834);
  and AND_9523(g14097,g878,g10632);
  and AND_9524(g14126,g881,g10632);
  and AND_9525(g14148,g884,g10632);
  and AND_9526(g14168,g887,g10632);
  and AND_9527(g14180,g872,g10632);
  and AND_9528(g14185,g8686,g11744);
  and AND_9529(g14190,g859,g10632);
  and AND_9530(g14193,g7178,g10590);
  and AND_9531(g14202,g869,g10632);
  and AND_9532(g14206,g8655,g11790);
  and AND_9533(g14207,g8639,g11793);
  and AND_9534(g14210,g4392,g10590);
  and AND_9535(g14216,g7631,g10608);
  and AND_9536(g14218,g875,g10632);
  and AND_9537(g14220,g8612,g11820);
  and AND_9538(g14221,g8686,g11823);
  and AND_9539(g14222,g8655,g11826);
  and AND_9540(g14233,g8639,g11855);
  and AND_9541(g14256,g2079,g11872);
  and AND_9542(g14257,g8612,g11878);
  and AND_9543(g14261,g4507,g10738);
  and AND_9544(g14295,g1811,g11894);
  and AND_9545(g14296,g2638,g11897);
  and AND_9546(g14316,g2370,g11920);
  and AND_9547(g14438,g1087,g10726);
  and AND_9548(I16618,g10124,g12341,g12293);
  and AND_9549(g14496,g12411,g12244,g12197,I16618);
  and AND_9550(g14506,g1430,g10755);
  and AND_9551(I16646,g10160,g12413,g12343);
  and AND_9552(g14528,g12459,g12306,g12245,I16646);
  and AND_9553(g14537,g10550,g10529);
  and AND_9554(I16671,g10185,g12461,g12415);
  and AND_9555(g14555,g12521,g12356,g12307,I16671);
  and AND_9556(g14565,g11934,g11952);
  and AND_9557(g14566,g10566,g10551);
  and AND_9558(g14567,g10568,g10552);
  and AND_9559(I16695,g10207,g12523,g12463);
  and AND_9560(g14581,g12587,g12428,g12357,I16695);
  and AND_9561(g14585,g1141,g10905);
  and AND_9562(g14586,g11953,g11970);
  and AND_9563(g14587,g10584,g10567);
  and AND_9564(g14588,g11957,g11974);
  and AND_9565(g14589,g10586,g10569);
  and AND_9566(I16721,g10224,g12589,g12525);
  and AND_9567(g14608,g12638,g12476,g12429,I16721);
  and AND_9568(g14610,g1484,g10935);
  and AND_9569(g14612,g11971,g11993);
  and AND_9570(g14613,g10602,g10585);
  and AND_9571(g14614,g11975,g11997);
  and AND_9572(g14615,g10604,g10587);
  and AND_9573(g14641,g11994,g12020);
  and AND_9574(g14643,g11998,g12023);
  and AND_9575(g14644,g10610,g10605);
  and AND_9576(g14654,g7178,g10476);
  and AND_9577(g14680,g12024,g12053);
  and AND_9578(g14681,g4392,g10476);
  and AND_9579(g14708,g74,g12369);
  and AND_9580(g14719,g4392,g10830);
  and AND_9581(g14791,g1146,g10909);
  and AND_9582(g14831,g1152,g10909);
  and AND_9583(g14832,g1489,g10939);
  and AND_9584(g14874,g1099,g10909);
  and AND_9585(g14875,g1495,g10939);
  and AND_9586(g14913,g1442,g10939);
  and AND_9587(g15075,g12850,g12955);
  and AND_9588(g15076,g2130,g12955);
  and AND_9589(g15077,g2138,g12955);
  and AND_9590(g15078,g10361,g12955);
  and AND_9591(g15079,g2151,g12955);
  and AND_9592(g15080,g12855,g12983);
  and AND_9593(g15081,g2689,g12983);
  and AND_9594(g15082,g2697,g12983);
  and AND_9595(g15083,g10362,g12983);
  and AND_9596(g15084,g2710,g12983);
  and AND_9597(g15103,g4180,g14454);
  and AND_9598(g15104,g6955,g14454);
  and AND_9599(g15105,g4235,g14454);
  and AND_9600(g15107,g4258,g14454);
  and AND_9601(g15108,g4264,g14454);
  and AND_9602(g15109,g4269,g14454);
  and AND_9603(g15110,g4245,g14454);
  and AND_9604(g15111,g4281,g14454);
  and AND_9605(g15112,g4284,g14454);
  and AND_9606(g15113,g4291,g14454);
  and AND_9607(g15114,g4239,g14454);
  and AND_9608(g15115,g2946,g14454);
  and AND_9609(g15116,g4297,g14454);
  and AND_9610(g15117,g4300,g14454);
  and AND_9611(g15118,g4253,g14454);
  and AND_9612(g15119,g4249,g14454);
  and AND_9613(g15507,g10970,g13305);
  and AND_9614(g15567,g392,g13312);
  and AND_9615(g15574,g4311,g13202);
  and AND_9616(g15589,g411,g13334);
  and AND_9617(g15590,g3139,g13530);
  and AND_9618(g15611,g471,g13437);
  and AND_9619(g15612,g3143,g13530);
  and AND_9620(g15613,g3490,g13555);
  and AND_9621(g15631,g168,g13437);
  and AND_9622(g15632,g3494,g13555);
  and AND_9623(g15633,g3841,g13584);
  and AND_9624(g15650,g8362,g13413);
  and AND_9625(g15651,g429,g13414);
  and AND_9626(g15652,g174,g13437);
  and AND_9627(g15653,g3119,g13530);
  and AND_9628(g15654,g3845,g13584);
  and AND_9629(g15672,g433,g13458);
  and AND_9630(g15673,g182,g13437);
  and AND_9631(g15678,g1094,g13846);
  and AND_9632(g15679,g3470,g13555);
  and AND_9633(g15693,g269,g13474);
  and AND_9634(g15694,g457,g13437);
  and AND_9635(g15699,g1437,g13861);
  and AND_9636(g15700,g3089,g13483);
  and AND_9637(g15701,g3821,g13584);
  and AND_9638(g15703,g452,g13437);
  and AND_9639(g15704,g3440,g13504);
  and AND_9640(g15706,g13296,g13484);
  and AND_9641(g15707,g4082,g13506);
  and AND_9642(g15711,g460,g13437);
  and AND_9643(g15712,g3791,g13521);
  and AND_9644(g15716,g468,g13437);
  and AND_9645(g15722,g464,g13437);
  and AND_9646(g15738,g1111,g13260);
  and AND_9647(g15745,g686,g13223);
  and AND_9648(g15749,g1454,g13273);
  and AND_9649(g15757,g3207,g14066);
  and AND_9650(g15779,g13909,g11214);
  and AND_9651(g15783,g3215,g14098);
  and AND_9652(g15784,g3235,g13977);
  and AND_9653(g15785,g3558,g14107);
  and AND_9654(g15786,g13940,g11233);
  and AND_9655(g15793,g3219,g13873);
  and AND_9656(g15794,g3239,g14008);
  and AND_9657(g15795,g3566,g14130);
  and AND_9658(g15796,g3586,g14015);
  and AND_9659(g15797,g3909,g14139);
  and AND_9660(g15804,g3223,g13889);
  and AND_9661(g15805,g3243,g14041);
  and AND_9662(g15807,g3570,g13898);
  and AND_9663(g15808,g3590,g14048);
  and AND_9664(g15809,g3917,g14154);
  and AND_9665(g15810,g3937,g14055);
  and AND_9666(g15812,g3227,g13915);
  and AND_9667(g15813,g3247,g14069);
  and AND_9668(g15814,g3574,g13920);
  and AND_9669(g15815,g3594,g14075);
  and AND_9670(g15817,g3921,g13929);
  and AND_9671(g15818,g3941,g14082);
  and AND_9672(g15819,g3251,g14101);
  and AND_9673(g15820,g3578,g13955);
  and AND_9674(g15821,g3598,g14110);
  and AND_9675(g15822,g3925,g13960);
  and AND_9676(g15823,g3945,g14116);
  and AND_9677(g15836,g3187,g14104);
  and AND_9678(g15837,g3255,g14127);
  and AND_9679(g15838,g3602,g14133);
  and AND_9680(g15839,g3929,g13990);
  and AND_9681(g15840,g3949,g14142);
  and AND_9682(g15841,g4273,g13868);
  and AND_9683(g15847,g3191,g14005);
  and AND_9684(g15848,g3259,g13892);
  and AND_9685(g15849,g3538,g14136);
  and AND_9686(g15850,g3606,g14151);
  and AND_9687(g15851,g3953,g14157);
  and AND_9688(g15852,g13820,g13223);
  and AND_9689(g15856,g9056,g14223);
  and AND_9690(g15857,g3199,g14038);
  and AND_9691(g15858,g3542,g14045);
  and AND_9692(g15859,g3610,g13923);
  and AND_9693(g15860,g3889,g14160);
  and AND_9694(g15861,g3957,g14170);
  and AND_9695(g15863,g13762,g13223);
  and AND_9696(g15870,g3231,g13948);
  and AND_9697(g15871,g3203,g13951);
  and AND_9698(g15872,g9095,g14234);
  and AND_9699(g15873,g3550,g14072);
  and AND_9700(g15874,g3893,g14079);
  and AND_9701(g15875,g3961,g13963);
  and AND_9702(g15876,g13512,g13223);
  and AND_9703(g15880,g3211,g13980);
  and AND_9704(g15881,g3582,g13983);
  and AND_9705(g15882,g3554,g13986);
  and AND_9706(g15883,g9180,g14258);
  and AND_9707(g15884,g3901,g14113);
  and AND_9708(g15902,g441,g13975);
  and AND_9709(g15903,g13796,g13223);
  and AND_9710(g15911,g3111,g13530);
  and AND_9711(g15912,g3562,g14018);
  and AND_9712(g15913,g3933,g14021);
  and AND_9713(g15914,g3905,g14024);
  and AND_9714(g15936,g475,g13999);
  and AND_9715(g15937,g11950,g14387);
  and AND_9716(g15966,g3462,g13555);
  and AND_9717(g15967,g3913,g14058);
  and AND_9718(g15978,g246,g14032);
  and AND_9719(g15995,g13314,g1157,g10666);
  and AND_9720(g16023,g3813,g13584);
  and AND_9721(g16025,g446,g14063);
  and AND_9722(g16026,g854,g14065);
  and AND_9723(g16047,g13322,g1500,g10699);
  and AND_9724(g16098,g5148,g14238);
  and AND_9725(g16122,g9491,g14291);
  and AND_9726(g16125,g5152,g14238);
  and AND_9727(g16126,g5495,g14262);
  and AND_9728(g16128,g14333,g14166);
  and AND_9729(g16160,g5499,g14262);
  and AND_9730(g16161,g5841,g14297);
  and AND_9731(g16163,g14254,g14179);
  and AND_9732(g16176,g14596,g11779);
  and AND_9733(g16177,g5128,g14238);
  and AND_9734(g16178,g5845,g14297);
  and AND_9735(g16179,g6187,g14321);
  and AND_9736(g16184,g9285,g14183);
  and AND_9737(g16185,g3263,g14011);
  and AND_9738(g16190,g14626,g11810);
  and AND_9739(g16191,g5475,g14262);
  and AND_9740(g16192,g6191,g14321);
  and AND_9741(g16193,g6533,g14348);
  and AND_9742(I17529,g13156,g11450,g6756);
  and AND_9743(g16194,g11547,g6782,g11640,I17529);
  and AND_9744(g16199,g3614,g14051);
  and AND_9745(g16202,g86,g14197);
  and AND_9746(g16203,g5821,g14297);
  and AND_9747(g16204,g6537,g14348);
  and AND_9748(I17542,g13156,g6767,g6756);
  and AND_9749(g16205,g11547,g6782,g11640,I17542);
  and AND_9750(g16207,g9839,g14204);
  and AND_9751(g16208,g3965,g14085);
  and AND_9752(g16211,g5445,g14215);
  and AND_9753(g16212,g6167,g14321);
  and AND_9754(I17552,g13156,g11450,g11498);
  and AND_9755(g16213,g6772,g6782,g11640,I17552);
  and AND_9756(g16221,g5791,g14231);
  and AND_9757(g16222,g6513,g14348);
  and AND_9758(g16224,g14583,g14232);
  and AND_9759(g16233,g6137,g14251);
  and AND_9760(I17575,g13156,g11450,g6756);
  and AND_9761(g16234,g6772,g6782,g11640,I17575);
  and AND_9762(g16243,g6483,g14275);
  and AND_9763(I17585,g14988,g11450,g11498);
  and AND_9764(g16244,g11547,g11592,g6789,I17585);
  and AND_9765(g16245,g14278,g14708);
  and AND_9766(g16279,g4512,g14424);
  and AND_9767(I17606,g14988,g11450,g6756);
  and AND_9768(g16283,g11547,g11592,g6789,I17606);
  and AND_9769(g16303,g4527,g12921);
  and AND_9770(g16324,g13657,g182);
  and AND_9771(g16422,g8216,g13627);
  and AND_9772(g16427,g5216,g14876);
  and AND_9773(g16474,g8280,g13666);
  and AND_9774(g16483,g5224,g14915);
  and AND_9775(g16484,g5244,g14755);
  and AND_9776(g16485,g5563,g14924);
  and AND_9777(I17692,g14988,g11450,g6756);
  and AND_9778(g16486,g6772,g11592,g6789,I17692);
  and AND_9779(g16513,g8345,g13708);
  and AND_9780(g16516,g5228,g14627);
  and AND_9781(g16517,g5248,g14797);
  and AND_9782(g16518,g5571,g14956);
  and AND_9783(g16519,g5591,g14804);
  and AND_9784(g16520,g5909,g14965);
  and AND_9785(g16531,g5232,g14656);
  and AND_9786(g16532,g5252,g14841);
  and AND_9787(g16534,g5575,g14665);
  and AND_9788(g16535,g5595,g14848);
  and AND_9789(g16536,g5917,g14996);
  and AND_9790(g16537,g5937,g14855);
  and AND_9791(g16538,g6255,g15005);
  and AND_9792(I17741,g14988,g11450,g11498);
  and AND_9793(g16539,g11547,g6782,g6789,I17741);
  and AND_9794(g16590,g5236,g14683);
  and AND_9795(g16591,g5256,g14879);
  and AND_9796(g16592,g5579,g14688);
  and AND_9797(g16593,g5599,g14885);
  and AND_9798(g16595,g5921,g14697);
  and AND_9799(g16596,g5941,g14892);
  and AND_9800(g16597,g6263,g15021);
  and AND_9801(g16598,g6283,g14899);
  and AND_9802(g16599,g6601,g15030);
  and AND_9803(g16610,g5260,g14918);
  and AND_9804(g16611,g5583,g14727);
  and AND_9805(g16612,g5603,g14927);
  and AND_9806(g16613,g5925,g14732);
  and AND_9807(g16614,g5945,g14933);
  and AND_9808(g16616,g6267,g14741);
  and AND_9809(g16617,g6287,g14940);
  and AND_9810(g16618,g6609,g15039);
  and AND_9811(g16619,g6629,g14947);
  and AND_9812(g16621,g8278,g13821);
  and AND_9813(g16633,g5196,g14921);
  and AND_9814(g16634,g5264,g14953);
  and AND_9815(g16635,g5607,g14959);
  and AND_9816(g16636,g5929,g14768);
  and AND_9817(g16637,g5949,g14968);
  and AND_9818(g16638,g6271,g14773);
  and AND_9819(g16639,g6291,g14974);
  and AND_9820(g16641,g6613,g14782);
  and AND_9821(g16642,g6633,g14981);
  and AND_9822(g16653,g8343,g13850);
  and AND_9823(g16662,g4552,g14753);
  and AND_9824(g16666,g5200,g14794);
  and AND_9825(g16667,g5268,g14659);
  and AND_9826(g16668,g5543,g14962);
  and AND_9827(g16669,g5611,g14993);
  and AND_9828(g16670,g5953,g14999);
  and AND_9829(g16671,g6275,g14817);
  and AND_9830(g16672,g6295,g15008);
  and AND_9831(g16673,g6617,g14822);
  and AND_9832(g16674,g6637,g15014);
  and AND_9833(g16690,g8399,g13867);
  and AND_9834(g16699,g7134,g12933);
  and AND_9835(g16700,g5208,g14838);
  and AND_9836(g16701,g5547,g14845);
  and AND_9837(g16702,g5615,g14691);
  and AND_9838(g16703,g5889,g15002);
  and AND_9839(g16704,g5957,g15018);
  and AND_9840(g16705,g6299,g15024);
  and AND_9841(g16706,g6621,g14868);
  and AND_9842(g16707,g6641,g15033);
  and AND_9843(g16729,g5240,g14720);
  and AND_9844(g16730,g5212,g14723);
  and AND_9845(g16731,g7153,g12941);
  and AND_9846(g16732,g5555,g14882);
  and AND_9847(g16733,g5893,g14889);
  and AND_9848(g16734,g5961,g14735);
  and AND_9849(g16735,g6235,g15027);
  and AND_9850(g16736,g6303,g15036);
  and AND_9851(g16737,g6645,g15042);
  and AND_9852(g16751,g13155,g13065);
  and AND_9853(g16758,g5220,g14758);
  and AND_9854(g16759,g5587,g14761);
  and AND_9855(g16760,g5559,g14764);
  and AND_9856(g16761,g7170,g12947);
  and AND_9857(g16762,g5901,g14930);
  and AND_9858(g16763,g6239,g14937);
  and AND_9859(g16764,g6307,g14776);
  and AND_9860(g16765,g6581,g15045);
  and AND_9861(g16766,g6649,g12915);
  and AND_9862(g16801,g5120,g14238);
  and AND_9863(g16802,g5567,g14807);
  and AND_9864(g16803,g5933,g14810);
  and AND_9865(g16804,g5905,g14813);
  and AND_9866(g16805,g7187,g12972);
  and AND_9867(g16806,g6247,g14971);
  and AND_9868(g16807,g6585,g14978);
  and AND_9869(g16808,g6653,g14825);
  and AND_9870(g16840,g5467,g14262);
  and AND_9871(g16841,g5913,g14858);
  and AND_9872(g16842,g6279,g14861);
  and AND_9873(g16843,g6251,g14864);
  and AND_9874(g16844,g7212,g13000);
  and AND_9875(g16845,g6593,g15011);
  and AND_9876(g16846,g14034,g12591,g11185);
  and AND_9877(g16855,g4392,g13107);
  and AND_9878(g16868,g5813,g14297);
  and AND_9879(g16869,g6259,g14902);
  and AND_9880(g16870,g6625,g14905);
  and AND_9881(g16871,g6597,g14908);
  and AND_9882(g16884,g6159,g14321);
  and AND_9883(g16885,g6605,g14950);
  and AND_9884(g16896,g262,g13120);
  and AND_9885(g16929,g6505,g14348);
  and AND_9886(g16930,g239,g13132);
  and AND_9887(g16957,g13064,g10418);
  and AND_9888(g16965,g269,g13140);
  and AND_9889(g16986,g246,g13142);
  and AND_9890(g17057,g446,g13173);
  and AND_9891(g17091,g8659,g12940);
  and AND_9892(g17119,g5272,g14800);
  and AND_9893(g17123,g225,g13209);
  and AND_9894(g17133,g10683,g13222);
  and AND_9895(g17134,g5619,g14851);
  and AND_9896(g17138,g255,g13239);
  and AND_9897(g17139,g8635,g12967);
  and AND_9898(g17140,g8616,g12968);
  and AND_9899(g17145,g7469,g13249);
  and AND_9900(g17146,g5965,g14895);
  and AND_9901(g17149,g232,g13255);
  and AND_9902(g17150,g8579,g12995);
  and AND_9903(g17151,g8659,g12996);
  and AND_9904(g17152,g8635,g12997);
  and AND_9905(g17153,g6311,g14943);
  and AND_9906(g17156,g305,g13385);
  and AND_9907(g17176,g8616,g13008);
  and AND_9908(g17177,g6657,g14984);
  and AND_9909(g17179,g1041,g13211);
  and AND_9910(g17181,g1945,g13014);
  and AND_9911(g17182,g8579,g13016);
  and AND_9912(g17191,g1384,g13242);
  and AND_9913(g17192,g1677,g13022);
  and AND_9914(g17193,g2504,g13023);
  and AND_9915(g17199,g2236,g13034);
  and AND_9916(g17292,g1075,g13093);
  and AND_9917(g17307,g9498,g14343);
  and AND_9918(g17317,g1079,g13124);
  and AND_9919(g17321,g1418,g13105);
  and AND_9920(g17365,g7650,g13036);
  and AND_9921(g17391,g9556,g14378);
  and AND_9922(g17401,g1083,g13143);
  and AND_9923(g17405,g1422,g13137);
  and AND_9924(g17418,g9618,g14407);
  and AND_9925(g17424,g1426,g13176);
  and AND_9926(g17469,g4076,g13217);
  and AND_9927(g17480,g9683,g14433);
  and AND_9928(g17506,g9744,g14505);
  and AND_9929(g17574,g9554,g14546);
  and AND_9930(g17601,g9616,g14572);
  and AND_9931(I18568,g13156,g11450,g11498);
  and AND_9932(g17613,g11547,g11592,g11640,I18568);
  and AND_9933(g17617,g7885,g13326);
  and AND_9934(g17636,g10829,g13463);
  and AND_9935(g17643,g9681,g14599);
  and AND_9936(I18620,g13156,g11450,g11498);
  and AND_9937(g17653,g11547,g11592,g6789,I18620);
  and AND_9938(g17654,g962,g13284);
  and AND_9939(g17655,g7897,g13342);
  and AND_9940(g17671,g7685,g13485);
  and AND_9941(g17682,g9742,g14637);
  and AND_9942(I18671,g13156,g11450,g6756);
  and AND_9943(g17690,g11547,g11592,g11640,I18671);
  and AND_9944(g17692,g1124,g13307);
  and AND_9945(g17693,g1306,g13291);
  and AND_9946(g17719,g9818,g14675);
  and AND_9947(I18713,g13156,g6767,g6756);
  and AND_9948(g17724,g11547,g11592,g11640,I18713);
  and AND_9949(I18716,g13156,g11450,g6756);
  and AND_9950(g17725,g11547,g11592,g6789,I18716);
  and AND_9951(g17726,g1467,g13315);
  and AND_9952(I18740,g13156,g11450,g11498);
  and AND_9953(g17747,g6772,g11592,g11640,I18740);
  and AND_9954(g17752,g7841,g13174);
  and AND_9955(g17753,g13281,g13175);
  and AND_9956(I18762,g13156,g6767,g11498);
  and AND_9957(g17766,g6772,g11592,g11640,I18762);
  and AND_9958(I18765,g13156,g11450,g11498);
  and AND_9959(g17767,g6772,g11592,g6789,I18765);
  and AND_9960(g17768,g13325,g10741);
  and AND_9961(g17769,g1146,g13188);
  and AND_9962(g17770,g7863,g13189);
  and AND_9963(g17771,g13288,g13190);
  and AND_9964(I18782,g13156,g11450,g6756);
  and AND_9965(g17780,g6772,g11592,g11640,I18782);
  and AND_9966(I18785,g13156,g6767,g11498);
  and AND_9967(g17781,g6772,g11592,g6789,I18785);
  and AND_9968(g17783,g7851,g13110);
  and AND_9969(g17784,g1152,g13215);
  and AND_9970(g17785,g13341,g10762);
  and AND_9971(g17786,g1489,g13216);
  and AND_9972(I18803,g13156,g11450,g6756);
  and AND_9973(g17793,g6772,g11592,g6789,I18803);
  and AND_9974(g17809,g7873,g13125);
  and AND_9975(g17810,g1495,g13246);
  and AND_9976(I18819,g13156,g11450,g11498);
  and AND_9977(g17817,g11547,g6782,g11640,I18819);
  and AND_9978(g18103,g401,g17015);
  and AND_9979(g18104,g392,g17015);
  and AND_9980(g18105,g417,g17015);
  and AND_9981(g18106,g411,g17015);
  and AND_9982(g18107,g429,g17015);
  and AND_9983(g18108,g433,g17015);
  and AND_9984(g18109,g437,g17015);
  and AND_9985(g18110,g441,g17015);
  and AND_9986(g18111,g174,g17015);
  and AND_9987(g18112,g182,g17015);
  and AND_9988(g18113,g405,g17015);
  and AND_9989(g18114,g452,g17015);
  and AND_9990(g18115,g460,g17015);
  and AND_9991(g18116,g168,g17015);
  and AND_9992(g18117,g464,g17015);
  and AND_9993(g18118,g471,g17015);
  and AND_9994(g18119,g475,g17015);
  and AND_9995(g18120,g457,g17015);
  and AND_9996(g18121,g424,g17015);
  and AND_9997(g18122,g15052,g17015);
  and AND_9998(g18123,g479,g16886);
  and AND_9999(g18124,g102,g16886);
  and AND_10000(g18125,g15053,g16886);
  and AND_10001(g18126,g15054,g16971);
  and AND_10002(g18127,g499,g16971);
  and AND_10003(g18128,g504,g16971);
  and AND_10004(g18129,g518,g16971);
  and AND_10005(g18130,g528,g16971);
  and AND_10006(g18131,g482,g16971);
  and AND_10007(g18132,g513,g16971);
  and AND_10008(g18133,g15055,g17249);
  and AND_10009(g18134,g534,g17249);
  and AND_10010(g18135,g136,g17249);
  and AND_10011(g18136,g550,g17249);
  and AND_10012(g18137,g538,g17249);
  and AND_10013(g18138,g546,g17249);
  and AND_10014(g18139,g542,g17249);
  and AND_10015(g18140,g559,g17533);
  and AND_10016(g18141,g568,g17533);
  and AND_10017(g18142,g577,g17533);
  and AND_10018(g18143,g586,g17533);
  and AND_10019(g18144,g590,g17533);
  and AND_10020(g18145,g582,g17533);
  and AND_10021(g18146,g595,g17533);
  and AND_10022(g18147,g599,g17533);
  and AND_10023(g18148,g562,g17533);
  and AND_10024(g18149,g608,g17533);
  and AND_10025(g18150,g604,g17533);
  and AND_10026(g18151,g617,g17533);
  and AND_10027(g18152,g613,g17533);
  and AND_10028(g18153,g626,g17533);
  and AND_10029(g18154,g622,g17533);
  and AND_10030(g18155,g15056,g17533);
  and AND_10031(g18156,g572,g17533);
  and AND_10032(g18157,g15057,g17433);
  and AND_10033(g18158,g667,g17433);
  and AND_10034(g18159,g671,g17433);
  and AND_10035(g18160,g645,g17433);
  and AND_10036(g18161,g691,g17433);
  and AND_10037(g18162,g686,g17433);
  and AND_10038(g18163,g79,g17433);
  and AND_10039(g18164,g699,g17433);
  and AND_10040(g18165,g650,g17433);
  and AND_10041(g18166,g655,g17433);
  and AND_10042(g18167,g718,g17433);
  and AND_10043(g18168,g681,g17433);
  and AND_10044(g18169,g676,g17433);
  and AND_10045(g18170,g661,g17433);
  and AND_10046(g18171,g728,g17433);
  and AND_10047(g18172,g15058,g17328);
  and AND_10048(g18173,g736,g17328);
  and AND_10049(g18174,g739,g17328);
  and AND_10050(g18175,g744,g17328);
  and AND_10051(g18176,g732,g17328);
  and AND_10052(g18177,g749,g17328);
  and AND_10053(g18178,g758,g17328);
  and AND_10054(g18179,g763,g17328);
  and AND_10055(g18180,g767,g17328);
  and AND_10056(g18181,g772,g17328);
  and AND_10057(g18182,g776,g17328);
  and AND_10058(g18183,g781,g17328);
  and AND_10059(g18184,g785,g17328);
  and AND_10060(g18185,g790,g17328);
  and AND_10061(g18186,g753,g17328);
  and AND_10062(g18187,g794,g17328);
  and AND_10063(g18188,g807,g17328);
  and AND_10064(g18189,g812,g17821);
  and AND_10065(g18190,g822,g17821);
  and AND_10066(g18191,g827,g17821);
  and AND_10067(g18192,g817,g17821);
  and AND_10068(g18193,g837,g17821);
  and AND_10069(g18194,g843,g17821);
  and AND_10070(g18195,g847,g17821);
  and AND_10071(g18196,g703,g17821);
  and AND_10072(g18197,g854,g17821);
  and AND_10073(g18198,g15059,g17821);
  and AND_10074(g18199,g832,g17821);
  and AND_10075(g18201,g15061,g15938);
  and AND_10076(g18202,g907,g15938);
  and AND_10077(g18203,g911,g15938);
  and AND_10078(g18204,g914,g15938);
  and AND_10079(g18205,g904,g15938);
  and AND_10080(g18206,g918,g15938);
  and AND_10081(g18207,g925,g15938);
  and AND_10082(g18208,g930,g15938);
  and AND_10083(g18209,g921,g15938);
  and AND_10084(g18210,g936,g15938);
  and AND_10085(g18211,g15062,g15979);
  and AND_10086(g18212,g947,g15979);
  and AND_10087(g18213,g952,g15979);
  and AND_10088(g18214,g939,g15979);
  and AND_10089(g18215,g943,g15979);
  and AND_10090(g18216,g967,g15979);
  and AND_10091(g18217,g15063,g16100);
  and AND_10092(g18218,g1008,g16100);
  and AND_10093(g18219,g969,g16100);
  and AND_10094(g18220,g1002,g16100);
  and AND_10095(g18221,g1018,g16100);
  and AND_10096(g18222,g1024,g16100);
  and AND_10097(g18223,g1030,g16100);
  and AND_10098(g18224,g1036,g16100);
  and AND_10099(g18225,g1041,g16100);
  and AND_10100(g18226,g15064,g16129);
  and AND_10101(g18227,g1052,g16129);
  and AND_10102(g18228,g1061,g16129);
  and AND_10103(g18229,g1099,g16326);
  and AND_10104(g18230,g1111,g16326);
  and AND_10105(g18231,g1105,g16326);
  and AND_10106(g18232,g1124,g16326);
  and AND_10107(g18233,g1094,g16326);
  and AND_10108(g18234,g1129,g16326);
  and AND_10109(g18235,g1141,g16326);
  and AND_10110(g18236,g15065,g16326);
  and AND_10111(g18237,g1146,g16326);
  and AND_10112(g18238,g1152,g16326);
  and AND_10113(g18239,g1135,g16326);
  and AND_10114(g18240,g15066,g16431);
  and AND_10115(g18241,g1183,g16431);
  and AND_10116(g18242,g962,g16431);
  and AND_10117(g18243,g1189,g16431);
  and AND_10118(g18244,g1171,g16431);
  and AND_10119(g18245,g1193,g16431);
  and AND_10120(g18246,g1199,g16431);
  and AND_10121(g18247,g1178,g16431);
  and AND_10122(g18248,g15067,g16897);
  and AND_10123(g18249,g1216,g16897);
  and AND_10124(g18250,g6821,g16897);
  and AND_10125(g18251,g996,g16897);
  and AND_10126(g18252,g990,g16897);
  and AND_10127(g18253,g1211,g16897);
  and AND_10128(g18254,g1236,g16897);
  and AND_10129(g18255,g1087,g16897);
  and AND_10130(g18256,g1242,g16897);
  and AND_10131(g18257,g1205,g16897);
  and AND_10132(g18258,g1221,g16897);
  and AND_10133(g18259,g15068,g16000);
  and AND_10134(g18260,g1252,g16000);
  and AND_10135(g18261,g1256,g16000);
  and AND_10136(g18262,g1259,g16000);
  and AND_10137(g18263,g1249,g16000);
  and AND_10138(g18264,g1263,g16000);
  and AND_10139(g18265,g1270,g16000);
  and AND_10140(g18266,g1274,g16000);
  and AND_10141(g18267,g1266,g16000);
  and AND_10142(g18268,g1280,g16000);
  and AND_10143(g18269,g15069,g16031);
  and AND_10144(g18270,g1291,g16031);
  and AND_10145(g18271,g1296,g16031);
  and AND_10146(g18272,g1283,g16031);
  and AND_10147(g18273,g1287,g16031);
  and AND_10148(g18274,g1311,g16031);
  and AND_10149(g18275,g15070,g16136);
  and AND_10150(g18276,g1351,g16136);
  and AND_10151(g18277,g1312,g16136);
  and AND_10152(g18278,g1345,g16136);
  and AND_10153(g18279,g1361,g16136);
  and AND_10154(g18280,g1367,g16136);
  and AND_10155(g18281,g1373,g16136);
  and AND_10156(g18282,g1379,g16136);
  and AND_10157(g18283,g1384,g16136);
  and AND_10158(g18284,g15071,g16164);
  and AND_10159(g18285,g1395,g16164);
  and AND_10160(g18286,g1404,g16164);
  and AND_10161(g18287,g1442,g16449);
  and AND_10162(g18288,g1454,g16449);
  and AND_10163(g18289,g1448,g16449);
  and AND_10164(g18290,g1467,g16449);
  and AND_10165(g18291,g1437,g16449);
  and AND_10166(g18292,g1472,g16449);
  and AND_10167(g18293,g1484,g16449);
  and AND_10168(g18294,g15072,g16449);
  and AND_10169(g18295,g1489,g16449);
  and AND_10170(g18296,g1495,g16449);
  and AND_10171(g18297,g1478,g16449);
  and AND_10172(g18298,g15073,g16489);
  and AND_10173(g18299,g1526,g16489);
  and AND_10174(g18300,g1306,g16489);
  and AND_10175(g18301,g1532,g16489);
  and AND_10176(g18302,g1514,g16489);
  and AND_10177(g18303,g1536,g16489);
  and AND_10178(g18304,g1542,g16489);
  and AND_10179(g18305,g1521,g16489);
  and AND_10180(g18306,g15074,g16931);
  and AND_10181(g18307,g1559,g16931);
  and AND_10182(g18308,g6832,g16931);
  and AND_10183(g18309,g1339,g16931);
  and AND_10184(g18310,g1333,g16931);
  and AND_10185(g18311,g1554,g16931);
  and AND_10186(g18312,g1579,g16931);
  and AND_10187(g18313,g1430,g16931);
  and AND_10188(g18314,g1585,g16931);
  and AND_10189(g18315,g1548,g16931);
  and AND_10190(g18316,g1564,g16931);
  and AND_10191(g18317,g12846,g17873);
  and AND_10192(g18318,g1604,g17873);
  and AND_10193(g18319,g1600,g17873);
  and AND_10194(g18320,g1616,g17873);
  and AND_10195(g18321,g1620,g17873);
  and AND_10196(g18322,g1608,g17873);
  and AND_10197(g18323,g1632,g17873);
  and AND_10198(g18324,g1644,g17873);
  and AND_10199(g18325,g1624,g17873);
  and AND_10200(g18326,g1664,g17873);
  and AND_10201(g18327,g1636,g17873);
  and AND_10202(g18328,g1657,g17873);
  and AND_10203(g18329,g1612,g17873);
  and AND_10204(g18330,g1668,g17873);
  and AND_10205(g18331,g1682,g17873);
  and AND_10206(g18332,g1677,g17873);
  and AND_10207(g18333,g1691,g17873);
  and AND_10208(g18334,g1696,g17873);
  and AND_10209(g18335,g1687,g17873);
  and AND_10210(g18336,g1700,g17873);
  and AND_10211(g18337,g1706,g17873);
  and AND_10212(g18338,g1710,g17873);
  and AND_10213(g18339,g1714,g17873);
  and AND_10214(g18340,g1720,g17873);
  and AND_10215(g18341,g1648,g17873);
  and AND_10216(g18342,g1592,g17873);
  and AND_10217(g18343,g12847,g17955);
  and AND_10218(g18344,g1740,g17955);
  and AND_10219(g18345,g1736,g17955);
  and AND_10220(g18346,g1752,g17955);
  and AND_10221(g18347,g1756,g17955);
  and AND_10222(g18348,g1744,g17955);
  and AND_10223(g18349,g1768,g17955);
  and AND_10224(g18350,g1779,g17955);
  and AND_10225(g18351,g1760,g17955);
  and AND_10226(g18352,g1798,g17955);
  and AND_10227(g18353,g1772,g17955);
  and AND_10228(g18354,g1792,g17955);
  and AND_10229(g18355,g1748,g17955);
  and AND_10230(g18356,g1802,g17955);
  and AND_10231(g18357,g1816,g17955);
  and AND_10232(g18358,g1811,g17955);
  and AND_10233(g18359,g1825,g17955);
  and AND_10234(g18360,g1830,g17955);
  and AND_10235(g18361,g1821,g17955);
  and AND_10236(g18362,g1834,g17955);
  and AND_10237(g18363,g1840,g17955);
  and AND_10238(g18364,g1844,g17955);
  and AND_10239(g18365,g1848,g17955);
  and AND_10240(g18366,g1854,g17955);
  and AND_10241(g18367,g1783,g17955);
  and AND_10242(g18368,g1728,g17955);
  and AND_10243(g18369,g12848,g15171);
  and AND_10244(g18370,g1874,g15171);
  and AND_10245(g18371,g1870,g15171);
  and AND_10246(g18372,g1886,g15171);
  and AND_10247(g18373,g1890,g15171);
  and AND_10248(g18374,g1878,g15171);
  and AND_10249(g18375,g1902,g15171);
  and AND_10250(g18376,g1913,g15171);
  and AND_10251(g18377,g1894,g15171);
  and AND_10252(g18378,g1932,g15171);
  and AND_10253(g18379,g1906,g15171);
  and AND_10254(g18380,g1926,g15171);
  and AND_10255(g18381,g1882,g15171);
  and AND_10256(g18382,g1936,g15171);
  and AND_10257(g18383,g1950,g15171);
  and AND_10258(g18384,g1945,g15171);
  and AND_10259(g18385,g1959,g15171);
  and AND_10260(g18386,g1964,g15171);
  and AND_10261(g18387,g1955,g15171);
  and AND_10262(g18388,g1968,g15171);
  and AND_10263(g18389,g1974,g15171);
  and AND_10264(g18390,g1978,g15171);
  and AND_10265(g18391,g1982,g15171);
  and AND_10266(g18392,g1988,g15171);
  and AND_10267(g18393,g1917,g15171);
  and AND_10268(g18394,g1862,g15171);
  and AND_10269(g18395,g12849,g15373);
  and AND_10270(g18396,g2008,g15373);
  and AND_10271(g18397,g2004,g15373);
  and AND_10272(g18398,g2020,g15373);
  and AND_10273(g18399,g2024,g15373);
  and AND_10274(g18400,g2012,g15373);
  and AND_10275(g18401,g2036,g15373);
  and AND_10276(g18402,g2047,g15373);
  and AND_10277(g18403,g2028,g15373);
  and AND_10278(g18404,g2066,g15373);
  and AND_10279(g18405,g2040,g15373);
  and AND_10280(g18406,g2060,g15373);
  and AND_10281(g18407,g2016,g15373);
  and AND_10282(g18408,g2070,g15373);
  and AND_10283(g18409,g2084,g15373);
  and AND_10284(g18410,g2079,g15373);
  and AND_10285(g18411,g2093,g15373);
  and AND_10286(g18412,g2098,g15373);
  and AND_10287(g18413,g2089,g15373);
  and AND_10288(g18414,g2102,g15373);
  and AND_10289(g18415,g2108,g15373);
  and AND_10290(g18416,g2112,g15373);
  and AND_10291(g18417,g2116,g15373);
  and AND_10292(g18418,g2122,g15373);
  and AND_10293(g18419,g2051,g15373);
  and AND_10294(g18420,g1996,g15373);
  and AND_10295(g18423,g12851,g18008);
  and AND_10296(g18424,g2165,g18008);
  and AND_10297(g18425,g2161,g18008);
  and AND_10298(g18426,g2177,g18008);
  and AND_10299(g18427,g2181,g18008);
  and AND_10300(g18428,g2169,g18008);
  and AND_10301(g18429,g2193,g18008);
  and AND_10302(g18430,g2204,g18008);
  and AND_10303(g18431,g2185,g18008);
  and AND_10304(g18432,g2223,g18008);
  and AND_10305(g18433,g2197,g18008);
  and AND_10306(g18434,g2217,g18008);
  and AND_10307(g18435,g2173,g18008);
  and AND_10308(g18436,g2227,g18008);
  and AND_10309(g18437,g2241,g18008);
  and AND_10310(g18438,g2236,g18008);
  and AND_10311(g18439,g2250,g18008);
  and AND_10312(g18440,g2255,g18008);
  and AND_10313(g18441,g2246,g18008);
  and AND_10314(g18442,g2259,g18008);
  and AND_10315(g18443,g2265,g18008);
  and AND_10316(g18444,g2269,g18008);
  and AND_10317(g18445,g2273,g18008);
  and AND_10318(g18446,g2279,g18008);
  and AND_10319(g18447,g2208,g18008);
  and AND_10320(g18448,g2153,g18008);
  and AND_10321(g18449,g12852,g15224);
  and AND_10322(g18450,g2299,g15224);
  and AND_10323(g18451,g2295,g15224);
  and AND_10324(g18452,g2311,g15224);
  and AND_10325(g18453,g2315,g15224);
  and AND_10326(g18454,g2303,g15224);
  and AND_10327(g18455,g2327,g15224);
  and AND_10328(g18456,g2338,g15224);
  and AND_10329(g18457,g2319,g15224);
  and AND_10330(g18458,g2357,g15224);
  and AND_10331(g18459,g2331,g15224);
  and AND_10332(g18460,g2351,g15224);
  and AND_10333(g18461,g2307,g15224);
  and AND_10334(g18462,g2361,g15224);
  and AND_10335(g18463,g2375,g15224);
  and AND_10336(g18464,g2370,g15224);
  and AND_10337(g18465,g2384,g15224);
  and AND_10338(g18466,g2389,g15224);
  and AND_10339(g18467,g2380,g15224);
  and AND_10340(g18468,g2393,g15224);
  and AND_10341(g18469,g2399,g15224);
  and AND_10342(g18470,g2403,g15224);
  and AND_10343(g18471,g2407,g15224);
  and AND_10344(g18472,g2413,g15224);
  and AND_10345(g18473,g2342,g15224);
  and AND_10346(g18474,g2287,g15224);
  and AND_10347(g18475,g12853,g15426);
  and AND_10348(g18476,g2433,g15426);
  and AND_10349(g18477,g2429,g15426);
  and AND_10350(g18478,g2445,g15426);
  and AND_10351(g18479,g2449,g15426);
  and AND_10352(g18480,g2437,g15426);
  and AND_10353(g18481,g2461,g15426);
  and AND_10354(g18482,g2472,g15426);
  and AND_10355(g18483,g2453,g15426);
  and AND_10356(g18484,g2491,g15426);
  and AND_10357(g18485,g2465,g15426);
  and AND_10358(g18486,g2485,g15426);
  and AND_10359(g18487,g2441,g15426);
  and AND_10360(g18488,g2495,g15426);
  and AND_10361(g18489,g2509,g15426);
  and AND_10362(g18490,g2504,g15426);
  and AND_10363(g18491,g2518,g15426);
  and AND_10364(g18492,g2523,g15426);
  and AND_10365(g18493,g2514,g15426);
  and AND_10366(g18494,g2527,g15426);
  and AND_10367(g18495,g2533,g15426);
  and AND_10368(g18496,g2537,g15426);
  and AND_10369(g18497,g2541,g15426);
  and AND_10370(g18498,g2547,g15426);
  and AND_10371(g18499,g2476,g15426);
  and AND_10372(g18500,g2421,g15426);
  and AND_10373(g18501,g12854,g15509);
  and AND_10374(g18502,g2567,g15509);
  and AND_10375(g18503,g2563,g15509);
  and AND_10376(g18504,g2579,g15509);
  and AND_10377(g18505,g2583,g15509);
  and AND_10378(g18506,g2571,g15509);
  and AND_10379(g18507,g2595,g15509);
  and AND_10380(g18508,g2606,g15509);
  and AND_10381(g18509,g2587,g15509);
  and AND_10382(g18510,g2625,g15509);
  and AND_10383(g18511,g2599,g15509);
  and AND_10384(g18512,g2619,g15509);
  and AND_10385(g18513,g2575,g15509);
  and AND_10386(g18514,g2629,g15509);
  and AND_10387(g18515,g2643,g15509);
  and AND_10388(g18516,g2638,g15509);
  and AND_10389(g18517,g2652,g15509);
  and AND_10390(g18518,g2657,g15509);
  and AND_10391(g18519,g2648,g15509);
  and AND_10392(g18520,g2661,g15509);
  and AND_10393(g18521,g2667,g15509);
  and AND_10394(g18522,g2671,g15509);
  and AND_10395(g18523,g2675,g15509);
  and AND_10396(g18524,g2681,g15509);
  and AND_10397(g18525,g2610,g15509);
  and AND_10398(g18526,g2555,g15509);
  and AND_10399(g18529,g2712,g15277);
  and AND_10400(g18530,g2715,g15277);
  and AND_10401(g18531,g2719,g15277);
  and AND_10402(g18532,g2724,g15277);
  and AND_10403(g18533,g2729,g15277);
  and AND_10404(g18534,g2735,g15277);
  and AND_10405(g18535,g2741,g15277);
  and AND_10406(g18536,g2748,g15277);
  and AND_10407(g18537,g6856,g15277);
  and AND_10408(g18538,g2759,g15277);
  and AND_10409(g18539,g2763,g15277);
  and AND_10410(g18540,g2775,g15277);
  and AND_10411(g18541,g2767,g15277);
  and AND_10412(g18542,g2787,g15277);
  and AND_10413(g18543,g2779,g15277);
  and AND_10414(g18544,g2791,g15277);
  and AND_10415(g18545,g2783,g15277);
  and AND_10416(g18546,g2795,g15277);
  and AND_10417(g18547,g121,g15277);
  and AND_10418(g18548,g2807,g15277);
  and AND_10419(g18549,g2799,g15277);
  and AND_10420(g18550,g2819,g15277);
  and AND_10421(g18551,g2811,g15277);
  and AND_10422(g18552,g2815,g15277);
  and AND_10423(g18553,g2827,g15277);
  and AND_10424(g18554,g2831,g15277);
  and AND_10425(g18555,g2834,g15277);
  and AND_10426(g18556,g2823,g15277);
  and AND_10427(g18557,g2771,g15277);
  and AND_10428(g18558,g2803,g15277);
  and AND_10429(g18559,g12856,g15277);
  and AND_10430(g18560,g2837,g15277);
  and AND_10431(g18561,g2841,g15277);
  and AND_10432(g18563,g2890,g16349);
  and AND_10433(g18564,g2844,g16349);
  and AND_10434(g18565,g2852,g16349);
  and AND_10435(g18566,g2860,g16349);
  and AND_10436(g18567,g2894,g16349);
  and AND_10437(g18568,g37,g16349);
  and AND_10438(g18569,g94,g16349);
  and AND_10439(g18570,g2848,g16349);
  and AND_10440(g18571,g2856,g16349);
  and AND_10441(g18572,g2864,g16349);
  and AND_10442(g18573,g2898,g16349);
  and AND_10443(g18574,g2882,g16349);
  and AND_10444(g18575,g2878,g16349);
  and AND_10445(g18576,g2868,g16349);
  and AND_10446(g18577,g2988,g16349);
  and AND_10447(g18578,g2873,g16349);
  and AND_10448(g18579,g2984,g16349);
  and AND_10449(g18580,g2907,g16349);
  and AND_10450(g18581,g2912,g16349);
  and AND_10451(g18582,g2922,g16349);
  and AND_10452(g18583,g2936,g16349);
  and AND_10453(g18584,g2950,g16349);
  and AND_10454(g18585,g2960,g16349);
  and AND_10455(g18586,g2886,g16349);
  and AND_10456(g18587,g2980,g16349);
  and AND_10457(g18588,g2970,g16349);
  and AND_10458(g18589,g2902,g16349);
  and AND_10459(g18590,g2917,g16349);
  and AND_10460(g18591,g2965,g16349);
  and AND_10461(g18592,g2994,g16349);
  and AND_10462(g18593,g2999,g16349);
  and AND_10463(g18594,g12858,g16349);
  and AND_10464(g18595,g2927,g16349);
  and AND_10465(g18596,g2941,g16349);
  and AND_10466(g18597,g2975,g16349);
  and AND_10467(g18598,g3003,g16349);
  and AND_10468(g18599,g2955,g16349);
  and AND_10469(g18600,g3111,g16987);
  and AND_10470(g18601,g3106,g16987);
  and AND_10471(g18602,g3115,g16987);
  and AND_10472(g18603,g3119,g16987);
  and AND_10473(g18604,g3125,g16987);
  and AND_10474(g18605,g3129,g16987);
  and AND_10475(g18606,g3133,g16987);
  and AND_10476(g18607,g3139,g16987);
  and AND_10477(g18608,g15087,g16987);
  and AND_10478(g18609,g3147,g16987);
  and AND_10479(g18610,g15088,g17059);
  and AND_10480(g18611,g15090,g17200);
  and AND_10481(g18612,g3329,g17200);
  and AND_10482(g18613,g3338,g17200);
  and AND_10483(g18614,g3343,g17200);
  and AND_10484(g18615,g3347,g17200);
  and AND_10485(g18616,g6875,g17200);
  and AND_10486(g18617,g3462,g17062);
  and AND_10487(g18618,g3457,g17062);
  and AND_10488(g18619,g3466,g17062);
  and AND_10489(g18620,g3470,g17062);
  and AND_10490(g18621,g3476,g17062);
  and AND_10491(g18622,g3480,g17062);
  and AND_10492(g18623,g3484,g17062);
  and AND_10493(g18624,g3490,g17062);
  and AND_10494(g18625,g15092,g17062);
  and AND_10495(g18626,g3498,g17062);
  and AND_10496(g18627,g15093,g17093);
  and AND_10497(g18628,g15095,g17226);
  and AND_10498(g18629,g3680,g17226);
  and AND_10499(g18630,g3689,g17226);
  and AND_10500(g18631,g3694,g17226);
  and AND_10501(g18632,g3698,g17226);
  and AND_10502(g18633,g6905,g17226);
  and AND_10503(g18634,g3813,g17096);
  and AND_10504(g18635,g3808,g17096);
  and AND_10505(g18636,g3817,g17096);
  and AND_10506(g18637,g3821,g17096);
  and AND_10507(g18638,g3827,g17096);
  and AND_10508(g18639,g3831,g17096);
  and AND_10509(g18640,g3835,g17096);
  and AND_10510(g18641,g3841,g17096);
  and AND_10511(g18642,g15097,g17096);
  and AND_10512(g18643,g3849,g17096);
  and AND_10513(g18644,g15098,g17125);
  and AND_10514(g18645,g15100,g17271);
  and AND_10515(g18646,g4031,g17271);
  and AND_10516(g18647,g4040,g17271);
  and AND_10517(g18648,g4045,g17271);
  and AND_10518(g18649,g4049,g17271);
  and AND_10519(g18650,g6928,g17271);
  and AND_10520(g18651,g15102,g16249);
  and AND_10521(g18652,g4172,g16249);
  and AND_10522(g18653,g4176,g16249);
  and AND_10523(g18654,g4146,g16249);
  and AND_10524(g18655,g15106,g14454);
  and AND_10525(g18656,g15120,g17128);
  and AND_10526(g18657,g4308,g17128);
  and AND_10527(g18658,g15121,g17183);
  and AND_10528(g18659,g4366,g17183);
  and AND_10529(g18662,g15126,g17367);
  and AND_10530(g18663,g4311,g17367);
  and AND_10531(g18664,g4332,g17367);
  and AND_10532(g18665,g4584,g17367);
  and AND_10533(g18666,g4593,g17367);
  and AND_10534(g18667,g4601,g17367);
  and AND_10535(g18668,g4322,g17367);
  and AND_10536(g18669,g4608,g17367);
  and AND_10537(g18670,g4621,g15758);
  and AND_10538(g18671,g4628,g15758);
  and AND_10539(g18672,g15127,g15758);
  and AND_10540(g18673,g4643,g15758);
  and AND_10541(g18674,g4340,g15758);
  and AND_10542(g18675,g4349,g15758);
  and AND_10543(g18676,g4358,g15758);
  and AND_10544(g18677,g4639,g15758);
  and AND_10545(g18678,g66,g15758);
  and AND_10546(g18679,g4633,g15758);
  and AND_10547(g18680,g15128,g15885);
  and AND_10548(g18681,g4653,g15885);
  and AND_10549(g18682,g4646,g15885);
  and AND_10550(g18683,g4674,g15885);
  and AND_10551(g18684,g4681,g15885);
  and AND_10552(g18685,g4688,g15885);
  and AND_10553(g18686,g4659,g15885);
  and AND_10554(g18687,g4664,g15885);
  and AND_10555(g18688,g4704,g16752);
  and AND_10556(g18689,g15129,g16752);
  and AND_10557(g18690,g15130,g16053);
  and AND_10558(g18691,g4727,g16053);
  and AND_10559(g18692,g4732,g16053);
  and AND_10560(g18693,g4717,g16053);
  and AND_10561(g18694,g4722,g16053);
  and AND_10562(g18695,g4737,g16053);
  and AND_10563(g18696,g4741,g16053);
  and AND_10564(g18697,g4749,g16777);
  and AND_10565(g18698,g15131,g16777);
  and AND_10566(g18699,g4760,g16816);
  and AND_10567(g18700,g15132,g16816);
  and AND_10568(g18701,g4771,g16856);
  and AND_10569(g18702,g15133,g16856);
  and AND_10570(g18703,g4776,g16782);
  and AND_10571(g18704,g4793,g16782);
  and AND_10572(g18705,g4801,g16782);
  and AND_10573(g18706,g4785,g16782);
  and AND_10574(g18707,g15134,g16782);
  and AND_10575(g18708,g4818,g16782);
  and AND_10576(g18709,g59,g17302);
  and AND_10577(g18710,g15135,g17302);
  and AND_10578(g18711,g15136,g15915);
  and AND_10579(g18712,g4843,g15915);
  and AND_10580(g18713,g4836,g15915);
  and AND_10581(g18714,g4864,g15915);
  and AND_10582(g18715,g4871,g15915);
  and AND_10583(g18716,g4878,g15915);
  and AND_10584(g18717,g4849,g15915);
  and AND_10585(g18718,g4854,g15915);
  and AND_10586(g18719,g4894,g16795);
  and AND_10587(g18720,g15137,g16795);
  and AND_10588(g18721,g15138,g16077);
  and AND_10589(g18722,g4917,g16077);
  and AND_10590(g18723,g4922,g16077);
  and AND_10591(g18724,g4907,g16077);
  and AND_10592(g18725,g4912,g16077);
  and AND_10593(g18726,g4927,g16077);
  and AND_10594(g18727,g4931,g16077);
  and AND_10595(g18728,g4939,g16821);
  and AND_10596(g18729,g15139,g16821);
  and AND_10597(g18730,g4950,g16861);
  and AND_10598(g18731,g15140,g16861);
  and AND_10599(g18732,g4961,g16877);
  and AND_10600(g18733,g15141,g16877);
  and AND_10601(g18734,g4966,g16826);
  and AND_10602(g18735,g4983,g16826);
  and AND_10603(g18736,g4991,g16826);
  and AND_10604(g18737,g4975,g16826);
  and AND_10605(g18738,g15142,g16826);
  and AND_10606(g18739,g5008,g16826);
  and AND_10607(g18740,g4572,g17384);
  and AND_10608(g18741,g15143,g17384);
  and AND_10609(g18742,g5120,g17847);
  and AND_10610(g18743,g5115,g17847);
  and AND_10611(g18744,g5124,g17847);
  and AND_10612(g18745,g5128,g17847);
  and AND_10613(g18746,g5134,g17847);
  and AND_10614(g18747,g5138,g17847);
  and AND_10615(g18748,g5142,g17847);
  and AND_10616(g18749,g5148,g17847);
  and AND_10617(g18750,g15145,g17847);
  and AND_10618(g18751,g5156,g17847);
  and AND_10619(g18752,g15146,g17926);
  and AND_10620(g18753,g15148,g15595);
  and AND_10621(g18754,g5339,g15595);
  and AND_10622(g18755,g5343,g15595);
  and AND_10623(g18756,g5348,g15595);
  and AND_10624(g18757,g5352,g15595);
  and AND_10625(g18758,g7004,g15595);
  and AND_10626(g18759,g5467,g17929);
  and AND_10627(g18760,g5462,g17929);
  and AND_10628(g18761,g5471,g17929);
  and AND_10629(g18762,g5475,g17929);
  and AND_10630(g18763,g5481,g17929);
  and AND_10631(g18764,g5485,g17929);
  and AND_10632(g18765,g5489,g17929);
  and AND_10633(g18766,g5495,g17929);
  and AND_10634(g18767,g15150,g17929);
  and AND_10635(g18768,g5503,g17929);
  and AND_10636(g18769,g15151,g18062);
  and AND_10637(g18770,g15153,g15615);
  and AND_10638(g18771,g5685,g15615);
  and AND_10639(g18772,g5689,g15615);
  and AND_10640(g18773,g5694,g15615);
  and AND_10641(g18774,g5698,g15615);
  and AND_10642(g18775,g7028,g15615);
  and AND_10643(g18776,g5813,g18065);
  and AND_10644(g18777,g5808,g18065);
  and AND_10645(g18778,g5817,g18065);
  and AND_10646(g18779,g5821,g18065);
  and AND_10647(g18780,g5827,g18065);
  and AND_10648(g18781,g5831,g18065);
  and AND_10649(g18782,g5835,g18065);
  and AND_10650(g18783,g5841,g18065);
  and AND_10651(g18784,g15155,g18065);
  and AND_10652(g18785,g5849,g18065);
  and AND_10653(g18786,g15156,g15345);
  and AND_10654(g18787,g15158,g15634);
  and AND_10655(g18788,g6031,g15634);
  and AND_10656(g18789,g6035,g15634);
  and AND_10657(g18790,g6040,g15634);
  and AND_10658(g18791,g6044,g15634);
  and AND_10659(g18792,g7051,g15634);
  and AND_10660(g18793,g6159,g15348);
  and AND_10661(g18794,g6154,g15348);
  and AND_10662(g18795,g6163,g15348);
  and AND_10663(g18796,g6167,g15348);
  and AND_10664(g18797,g6173,g15348);
  and AND_10665(g18798,g6177,g15348);
  and AND_10666(g18799,g6181,g15348);
  and AND_10667(g18800,g6187,g15348);
  and AND_10668(g18801,g15160,g15348);
  and AND_10669(g18802,g6195,g15348);
  and AND_10670(g18803,g15161,g15480);
  and AND_10671(g18804,g15163,g15656);
  and AND_10672(g18805,g6377,g15656);
  and AND_10673(g18806,g6381,g15656);
  and AND_10674(g18807,g6386,g15656);
  and AND_10675(g18808,g6390,g15656);
  and AND_10676(g18809,g7074,g15656);
  and AND_10677(g18810,g6505,g15483);
  and AND_10678(g18811,g6500,g15483);
  and AND_10679(g18812,g6509,g15483);
  and AND_10680(g18813,g6513,g15483);
  and AND_10681(g18814,g6519,g15483);
  and AND_10682(g18815,g6523,g15483);
  and AND_10683(g18816,g6527,g15483);
  and AND_10684(g18817,g6533,g15483);
  and AND_10685(g18818,g15165,g15483);
  and AND_10686(g18819,g6541,g15483);
  and AND_10687(g18820,g15166,g15563);
  and AND_10688(g18821,g15168,g15680);
  and AND_10689(g18822,g6723,g15680);
  and AND_10690(g18823,g6727,g15680);
  and AND_10691(g18824,g6732,g15680);
  and AND_10692(g18825,g6736,g15680);
  and AND_10693(g18826,g7097,g15680);
  and AND_10694(g18890,g10158,g17625);
  and AND_10695(g18893,g16215,g16030);
  and AND_10696(g18906,g13568,g16264);
  and AND_10697(g18909,g16226,g13570);
  and AND_10698(g18910,g16227,g16075);
  and AND_10699(g18933,g16237,g13597);
  and AND_10700(g18934,g3133,g16096);
  and AND_10701(g18935,g4322,g15574);
  and AND_10702(g18943,g269,g16099);
  and AND_10703(g18949,g10183,g17625);
  and AND_10704(g18950,g11193,g16123);
  and AND_10705(g18951,g3484,g16124);
  and AND_10706(g18974,g174,g16127);
  and AND_10707(g18981,g11206,g16158);
  and AND_10708(g18982,g3835,g16159);
  and AND_10709(g18987,g182,g16162);
  and AND_10710(g18992,g8341,g16171);
  and AND_10711(g18993,g11224,g16172);
  and AND_10712(g19062,g446,g16180);
  and AND_10713(g19069,g8397,g16186);
  and AND_10714(g19139,g452,g16195);
  and AND_10715(g19145,g8450,g16200);
  and AND_10716(g19206,g460,g16206);
  and AND_10717(g19207,g7803,g15992);
  and AND_10718(g19266,g246,g16214);
  and AND_10719(g19275,g7823,g16044);
  and AND_10720(g19333,g464,g16223);
  and AND_10721(g19350,g15968,g13505);
  and AND_10722(g19354,g471,g16235);
  and AND_10723(g19372,g686,g16289);
  and AND_10724(g19383,g16893,g13223);
  and AND_10725(g19384,g667,g16310);
  and AND_10726(g19393,g691,g16325);
  and AND_10727(g19461,g11708,g16846);
  and AND_10728(g19462,g7850,g14182,g14177,g16646);
  and AND_10729(g19487,g499,g16680);
  and AND_10730(g19500,g504,g16712);
  and AND_10731(g19516,g7824,g16097);
  and AND_10732(g19521,g513,g16739);
  and AND_10733(g19536,g518,g16768);
  and AND_10734(g19540,g1124,g15904);
  and AND_10735(g19545,g3147,g16769);
  and AND_10736(g19556,g11932,g16809);
  and AND_10737(g19560,g15832,g1157,g10893);
  and AND_10738(g19564,g17175,g13976);
  and AND_10739(g19568,g1467,g15959);
  and AND_10740(g19571,g3498,g16812);
  and AND_10741(g19578,g16183,g11130);
  and AND_10742(g19581,g15843,g1500,g10918);
  and AND_10743(g19585,g17180,g14004);
  and AND_10744(g19588,g3849,g16853);
  and AND_10745(g19594,g11913,g17268);
  and AND_10746(g19596,g1094,g16681);
  and AND_10747(g19601,g16198,g11149);
  and AND_10748(g19610,g1141,g16069);
  and AND_10749(g19613,g1437,g16713);
  and AND_10750(g19631,g1484,g16093);
  and AND_10751(g19637,g5142,g16958);
  and AND_10752(g19651,g1111,g16119);
  and AND_10753(g19655,g2729,g16966);
  and AND_10754(g19656,g2807,g15844);
  and AND_10755(g19660,g12001,g16968);
  and AND_10756(g19661,g5489,g16969);
  and AND_10757(g19671,g1454,g16155);
  and AND_10758(g19674,g2819,g15867);
  and AND_10759(g19680,g12028,g17013);
  and AND_10760(g19681,g5835,g17014);
  and AND_10761(g19684,g2735,g17297);
  and AND_10762(g19691,g9614,g17085);
  and AND_10763(g19692,g12066,g17086);
  and AND_10764(g19693,g6181,g17087);
  and AND_10765(g19715,g9679,g17120);
  and AND_10766(g19716,g12100,g17121);
  and AND_10767(g19717,g6527,g17122);
  and AND_10768(g19735,g9740,g17135);
  and AND_10769(g19736,g12136,g17136);
  and AND_10770(g19740,g2783,g15907);
  and AND_10771(g19746,g9816,g17147);
  and AND_10772(g19749,g732,g16646);
  and AND_10773(g19752,g2771,g15864);
  and AND_10774(g19756,g9899,g17154);
  and AND_10775(g19767,g16810,g14203);
  and AND_10776(g19768,g2803,g15833);
  and AND_10777(g19784,g2775,g15877);
  and AND_10778(g19788,g9983,g17216);
  and AND_10779(g19791,g14253,g17189);
  and AND_10780(g19855,g2787,g15962);
  and AND_10781(g19911,g14707,g17748);
  and AND_10782(g19914,g2815,g15853);
  and AND_10783(g19948,g17515,g16320);
  and AND_10784(g20056,g16291,g9007,g8954,g8903);
  and AND_10785(g20069,g16312,g9051,g9011,g8955);
  and AND_10786(g20084,g11591,g16609);
  and AND_10787(g20093,g15372,g14584);
  and AND_10788(g20094,g8872,g16631);
  and AND_10789(g20095,g8873,g16632);
  and AND_10790(g20108,g15508,g11048);
  and AND_10791(g20109,g17954,g17616);
  and AND_10792(g20112,g13540,g16661);
  and AND_10793(g20131,g15170,g14309);
  and AND_10794(g20135,g16258,g16695);
  and AND_10795(g20152,g11545,g16727);
  and AND_10796(g20162,g8737,g16750);
  and AND_10797(g20165,g5156,g17733);
  and AND_10798(g20171,g16479,g10476);
  and AND_10799(g20174,g5503,g17754);
  and AND_10800(g20188,g5849,g17772);
  and AND_10801(g20193,g15578,g17264);
  and AND_10802(g20203,g6195,g17789);
  and AND_10803(g20215,g16479,g10476);
  and AND_10804(g20218,g6541,g17815);
  and AND_10805(g20375,g671,g16846);
  and AND_10806(g20559,g336,g15831);
  and AND_10807(g20581,g10801,g15571);
  and AND_10808(g20602,g10803,g15580);
  and AND_10809(g20628,g1046,g15789);
  and AND_10810(g20658,g1389,g15800);
  and AND_10811(g20682,g16238,g4646);
  and AND_10812(g20739,g16259,g4674);
  and AND_10813(g20751,g16260,g4836);
  and AND_10814(g20875,g16281,g4681);
  and AND_10815(g20887,g16282,g4864);
  and AND_10816(g20977,g10123,g17301);
  and AND_10817(g21012,g16304,g4688);
  and AND_10818(g21024,g16306,g4871);
  and AND_10819(g21066,g10043,g17625);
  and AND_10820(g21067,g10085,g17625);
  and AND_10821(g21163,g16321,g4878);
  and AND_10822(g21188,g7666,g15705);
  and AND_10823(g21251,g13969,g17470);
  and AND_10824(g21276,g10157,g17625);
  and AND_10825(g21285,g7857,g16027);
  and AND_10826(g21296,g7879,g16072);
  and AND_10827(g21298,g7697,g15825);
  and AND_10828(g21302,g956,g15731);
  and AND_10829(g21303,g10120,g17625);
  and AND_10830(g21332,g996,g15739);
  and AND_10831(g21333,g1300,g15740);
  and AND_10832(g21347,g1339,g15750);
  and AND_10833(g21348,g10121,g17625);
  and AND_10834(g21361,g7869,g16066);
  and AND_10835(g21378,g7887,g16090);
  and AND_10836(g21382,g10086,g17625);
  and AND_10837(g21394,g13335,g15799);
  and AND_10838(g21404,g16069,g13569);
  and AND_10839(g21405,g13377,g15811);
  and AND_10840(g21419,g16681,g13595);
  and AND_10841(g21420,g16093,g13596);
  and AND_10842(g21452,g16119,g13624);
  and AND_10843(g21453,g16713,g13625);
  and AND_10844(g21464,g16181,g10872);
  and AND_10845(g21465,g16155,g13663);
  and AND_10846(g21512,g16225,g10881);
  and AND_10847(g21513,g16196,g10882);
  and AND_10848(g21557,g12980,g15674);
  and AND_10849(g21558,g15904,g13729);
  and AND_10850(g21559,g16236,g10897);
  and AND_10851(g21605,g13005,g15695);
  and AND_10852(g21606,g15959,g13763);
  and AND_10853(g21699,g142,g20283);
  and AND_10854(g21700,g150,g20283);
  and AND_10855(g21701,g153,g20283);
  and AND_10856(g21702,g157,g20283);
  and AND_10857(g21703,g146,g20283);
  and AND_10858(g21704,g164,g20283);
  and AND_10859(g21705,g209,g20283);
  and AND_10860(g21706,g222,g20283);
  and AND_10861(g21707,g191,g20283);
  and AND_10862(g21708,g15049,g20283);
  and AND_10863(g21709,g283,g20283);
  and AND_10864(g21710,g287,g20283);
  and AND_10865(g21711,g291,g20283);
  and AND_10866(g21712,g294,g20283);
  and AND_10867(g21713,g298,g20283);
  and AND_10868(g21714,g278,g20283);
  and AND_10869(g21715,g160,g20283);
  and AND_10870(g21716,g301,g20283);
  and AND_10871(g21717,g15051,g21037);
  and AND_10872(g21718,g370,g21037);
  and AND_10873(g21719,g358,g21037);
  and AND_10874(g21720,g376,g21037);
  and AND_10875(g21721,g385,g21037);
  and AND_10876(g21728,g3010,g20330);
  and AND_10877(g21729,g3021,g20330);
  and AND_10878(g21730,g3025,g20330);
  and AND_10879(g21731,g3029,g20330);
  and AND_10880(g21732,g3004,g20330);
  and AND_10881(g21733,g3034,g20330);
  and AND_10882(g21734,g3040,g20330);
  and AND_10883(g21735,g3057,g20330);
  and AND_10884(g21736,g3065,g20330);
  and AND_10885(g21737,g3068,g20330);
  and AND_10886(g21738,g3072,g20330);
  and AND_10887(g21739,g3080,g20330);
  and AND_10888(g21740,g3085,g20330);
  and AND_10889(g21741,g15086,g20330);
  and AND_10890(g21742,g3050,g20330);
  and AND_10891(g21743,g3100,g20330);
  and AND_10892(g21744,g3103,g20330);
  and AND_10893(g21745,g3017,g20330);
  and AND_10894(g21746,g3045,g20330);
  and AND_10895(g21747,g3061,g20330);
  and AND_10896(g21748,g15089,g20785);
  and AND_10897(g21749,g3155,g20785);
  and AND_10898(g21750,g3161,g20785);
  and AND_10899(g21751,g3167,g20785);
  and AND_10900(g21752,g3171,g20785);
  and AND_10901(g21753,g3179,g20785);
  and AND_10902(g21754,g3195,g20785);
  and AND_10903(g21755,g3203,g20785);
  and AND_10904(g21756,g3211,g20785);
  and AND_10905(g21757,g3187,g20785);
  and AND_10906(g21758,g3191,g20785);
  and AND_10907(g21759,g3199,g20785);
  and AND_10908(g21760,g3207,g20785);
  and AND_10909(g21761,g3215,g20785);
  and AND_10910(g21762,g3219,g20785);
  and AND_10911(g21763,g3223,g20785);
  and AND_10912(g21764,g3227,g20785);
  and AND_10913(g21765,g3231,g20785);
  and AND_10914(g21766,g3235,g20785);
  and AND_10915(g21767,g3239,g20785);
  and AND_10916(g21768,g3243,g20785);
  and AND_10917(g21769,g3247,g20785);
  and AND_10918(g21770,g3251,g20785);
  and AND_10919(g21771,g3255,g20785);
  and AND_10920(g21772,g3259,g20785);
  and AND_10921(g21773,g3263,g20785);
  and AND_10922(g21774,g3361,g20391);
  and AND_10923(g21775,g3372,g20391);
  and AND_10924(g21776,g3376,g20391);
  and AND_10925(g21777,g3380,g20391);
  and AND_10926(g21778,g3355,g20391);
  and AND_10927(g21779,g3385,g20391);
  and AND_10928(g21780,g3391,g20391);
  and AND_10929(g21781,g3408,g20391);
  and AND_10930(g21782,g3416,g20391);
  and AND_10931(g21783,g3419,g20391);
  and AND_10932(g21784,g3423,g20391);
  and AND_10933(g21785,g3431,g20391);
  and AND_10934(g21786,g3436,g20391);
  and AND_10935(g21787,g15091,g20391);
  and AND_10936(g21788,g3401,g20391);
  and AND_10937(g21789,g3451,g20391);
  and AND_10938(g21790,g3454,g20391);
  and AND_10939(g21791,g3368,g20391);
  and AND_10940(g21792,g3396,g20391);
  and AND_10941(g21793,g3412,g20391);
  and AND_10942(g21794,g15094,g20924);
  and AND_10943(g21795,g3506,g20924);
  and AND_10944(g21796,g3512,g20924);
  and AND_10945(g21797,g3518,g20924);
  and AND_10946(g21798,g3522,g20924);
  and AND_10947(g21799,g3530,g20924);
  and AND_10948(g21800,g3546,g20924);
  and AND_10949(g21801,g3554,g20924);
  and AND_10950(g21802,g3562,g20924);
  and AND_10951(g21803,g3538,g20924);
  and AND_10952(g21804,g3542,g20924);
  and AND_10953(g21805,g3550,g20924);
  and AND_10954(g21806,g3558,g20924);
  and AND_10955(g21807,g3566,g20924);
  and AND_10956(g21808,g3570,g20924);
  and AND_10957(g21809,g3574,g20924);
  and AND_10958(g21810,g3578,g20924);
  and AND_10959(g21811,g3582,g20924);
  and AND_10960(g21812,g3586,g20924);
  and AND_10961(g21813,g3590,g20924);
  and AND_10962(g21814,g3594,g20924);
  and AND_10963(g21815,g3598,g20924);
  and AND_10964(g21816,g3602,g20924);
  and AND_10965(g21817,g3606,g20924);
  and AND_10966(g21818,g3610,g20924);
  and AND_10967(g21819,g3614,g20924);
  and AND_10968(g21820,g3712,g20453);
  and AND_10969(g21821,g3723,g20453);
  and AND_10970(g21822,g3727,g20453);
  and AND_10971(g21823,g3731,g20453);
  and AND_10972(g21824,g3706,g20453);
  and AND_10973(g21825,g3736,g20453);
  and AND_10974(g21826,g3742,g20453);
  and AND_10975(g21827,g3759,g20453);
  and AND_10976(g21828,g3767,g20453);
  and AND_10977(g21829,g3770,g20453);
  and AND_10978(g21830,g3774,g20453);
  and AND_10979(g21831,g3782,g20453);
  and AND_10980(g21832,g3787,g20453);
  and AND_10981(g21833,g15096,g20453);
  and AND_10982(g21834,g3752,g20453);
  and AND_10983(g21835,g3802,g20453);
  and AND_10984(g21836,g3805,g20453);
  and AND_10985(g21837,g3719,g20453);
  and AND_10986(g21838,g3747,g20453);
  and AND_10987(g21839,g3763,g20453);
  and AND_10988(g21840,g15099,g21070);
  and AND_10989(g21841,g3857,g21070);
  and AND_10990(g21842,g3863,g21070);
  and AND_10991(g21843,g3869,g21070);
  and AND_10992(g21844,g3873,g21070);
  and AND_10993(g21845,g3881,g21070);
  and AND_10994(g21846,g3897,g21070);
  and AND_10995(g21847,g3905,g21070);
  and AND_10996(g21848,g3913,g21070);
  and AND_10997(g21849,g3889,g21070);
  and AND_10998(g21850,g3893,g21070);
  and AND_10999(g21851,g3901,g21070);
  and AND_11000(g21852,g3909,g21070);
  and AND_11001(g21853,g3917,g21070);
  and AND_11002(g21854,g3921,g21070);
  and AND_11003(g21855,g3925,g21070);
  and AND_11004(g21856,g3929,g21070);
  and AND_11005(g21857,g3933,g21070);
  and AND_11006(g21858,g3937,g21070);
  and AND_11007(g21859,g3941,g21070);
  and AND_11008(g21860,g3945,g21070);
  and AND_11009(g21861,g3949,g21070);
  and AND_11010(g21862,g3953,g21070);
  and AND_11011(g21863,g3957,g21070);
  and AND_11012(g21864,g3961,g21070);
  and AND_11013(g21865,g3965,g21070);
  and AND_11014(g21866,g4072,g19801);
  and AND_11015(g21867,g4082,g19801);
  and AND_11016(g21868,g4076,g19801);
  and AND_11017(g21869,g4087,g19801);
  and AND_11018(g21870,g4093,g19801);
  and AND_11019(g21871,g4108,g19801);
  and AND_11020(g21872,g4098,g19801);
  and AND_11021(g21873,g6946,g19801);
  and AND_11022(g21874,g4112,g19801);
  and AND_11023(g21875,g4116,g19801);
  and AND_11024(g21876,g4119,g19801);
  and AND_11025(g21877,g6888,g19801);
  and AND_11026(g21878,g4129,g19801);
  and AND_11027(g21879,g4132,g19801);
  and AND_11028(g21880,g4135,g19801);
  and AND_11029(g21881,g4064,g19801);
  and AND_11030(g21882,g4057,g19801);
  and AND_11031(g21883,g4141,g19801);
  and AND_11032(g21884,g4104,g19801);
  and AND_11033(g21885,g4122,g19801);
  and AND_11034(g21886,g4153,g19801);
  and AND_11035(g21887,g15101,g19801);
  and AND_11036(g21888,g4165,g19801);
  and AND_11037(g21889,g4169,g19801);
  and AND_11038(g21890,g4125,g19801);
  and AND_11039(g21906,g5022,g21468);
  and AND_11040(g21907,g5033,g21468);
  and AND_11041(g21908,g5037,g21468);
  and AND_11042(g21909,g5041,g21468);
  and AND_11043(g21910,g5016,g21468);
  and AND_11044(g21911,g5046,g21468);
  and AND_11045(g21912,g5052,g21468);
  and AND_11046(g21913,g5069,g21468);
  and AND_11047(g21914,g5077,g21468);
  and AND_11048(g21915,g5080,g21468);
  and AND_11049(g21916,g5084,g21468);
  and AND_11050(g21917,g5092,g21468);
  and AND_11051(g21918,g5097,g21468);
  and AND_11052(g21919,g15144,g21468);
  and AND_11053(g21920,g5062,g21468);
  and AND_11054(g21921,g5109,g21468);
  and AND_11055(g21922,g5112,g21468);
  and AND_11056(g21923,g5029,g21468);
  and AND_11057(g21924,g5057,g21468);
  and AND_11058(g21925,g5073,g21468);
  and AND_11059(g21926,g15147,g18997);
  and AND_11060(g21927,g5164,g18997);
  and AND_11061(g21928,g5170,g18997);
  and AND_11062(g21929,g5176,g18997);
  and AND_11063(g21930,g5180,g18997);
  and AND_11064(g21931,g5188,g18997);
  and AND_11065(g21932,g5204,g18997);
  and AND_11066(g21933,g5212,g18997);
  and AND_11067(g21934,g5220,g18997);
  and AND_11068(g21935,g5196,g18997);
  and AND_11069(g21936,g5200,g18997);
  and AND_11070(g21937,g5208,g18997);
  and AND_11071(g21938,g5216,g18997);
  and AND_11072(g21939,g5224,g18997);
  and AND_11073(g21940,g5228,g18997);
  and AND_11074(g21941,g5232,g18997);
  and AND_11075(g21942,g5236,g18997);
  and AND_11076(g21943,g5240,g18997);
  and AND_11077(g21944,g5244,g18997);
  and AND_11078(g21945,g5248,g18997);
  and AND_11079(g21946,g5252,g18997);
  and AND_11080(g21947,g5256,g18997);
  and AND_11081(g21948,g5260,g18997);
  and AND_11082(g21949,g5264,g18997);
  and AND_11083(g21950,g5268,g18997);
  and AND_11084(g21951,g5272,g18997);
  and AND_11085(g21952,g5366,g21514);
  and AND_11086(g21953,g5377,g21514);
  and AND_11087(g21954,g5381,g21514);
  and AND_11088(g21955,g5385,g21514);
  and AND_11089(g21956,g5360,g21514);
  and AND_11090(g21957,g5390,g21514);
  and AND_11091(g21958,g5396,g21514);
  and AND_11092(g21959,g5413,g21514);
  and AND_11093(g21960,g5421,g21514);
  and AND_11094(g21961,g5424,g21514);
  and AND_11095(g21962,g5428,g21514);
  and AND_11096(g21963,g5436,g21514);
  and AND_11097(g21964,g5441,g21514);
  and AND_11098(g21965,g15149,g21514);
  and AND_11099(g21966,g5406,g21514);
  and AND_11100(g21967,g5456,g21514);
  and AND_11101(g21968,g5459,g21514);
  and AND_11102(g21969,g5373,g21514);
  and AND_11103(g21970,g5401,g21514);
  and AND_11104(g21971,g5417,g21514);
  and AND_11105(g21972,g15152,g19074);
  and AND_11106(g21973,g5511,g19074);
  and AND_11107(g21974,g5517,g19074);
  and AND_11108(g21975,g5523,g19074);
  and AND_11109(g21976,g5527,g19074);
  and AND_11110(g21977,g5535,g19074);
  and AND_11111(g21978,g5551,g19074);
  and AND_11112(g21979,g5559,g19074);
  and AND_11113(g21980,g5567,g19074);
  and AND_11114(g21981,g5543,g19074);
  and AND_11115(g21982,g5547,g19074);
  and AND_11116(g21983,g5555,g19074);
  and AND_11117(g21984,g5563,g19074);
  and AND_11118(g21985,g5571,g19074);
  and AND_11119(g21986,g5575,g19074);
  and AND_11120(g21987,g5579,g19074);
  and AND_11121(g21988,g5583,g19074);
  and AND_11122(g21989,g5587,g19074);
  and AND_11123(g21990,g5591,g19074);
  and AND_11124(g21991,g5595,g19074);
  and AND_11125(g21992,g5599,g19074);
  and AND_11126(g21993,g5603,g19074);
  and AND_11127(g21994,g5607,g19074);
  and AND_11128(g21995,g5611,g19074);
  and AND_11129(g21996,g5615,g19074);
  and AND_11130(g21997,g5619,g19074);
  and AND_11131(g21998,g5712,g21562);
  and AND_11132(g21999,g5723,g21562);
  and AND_11133(g22000,g5727,g21562);
  and AND_11134(g22001,g5731,g21562);
  and AND_11135(g22002,g5706,g21562);
  and AND_11136(g22003,g5736,g21562);
  and AND_11137(g22004,g5742,g21562);
  and AND_11138(g22005,g5759,g21562);
  and AND_11139(g22006,g5767,g21562);
  and AND_11140(g22007,g5770,g21562);
  and AND_11141(g22008,g5774,g21562);
  and AND_11142(g22009,g5782,g21562);
  and AND_11143(g22010,g5787,g21562);
  and AND_11144(g22011,g15154,g21562);
  and AND_11145(g22012,g5752,g21562);
  and AND_11146(g22013,g5802,g21562);
  and AND_11147(g22014,g5805,g21562);
  and AND_11148(g22015,g5719,g21562);
  and AND_11149(g22016,g5747,g21562);
  and AND_11150(g22017,g5763,g21562);
  and AND_11151(g22018,g15157,g19147);
  and AND_11152(g22019,g5857,g19147);
  and AND_11153(g22020,g5863,g19147);
  and AND_11154(g22021,g5869,g19147);
  and AND_11155(g22022,g5873,g19147);
  and AND_11156(g22023,g5881,g19147);
  and AND_11157(g22024,g5897,g19147);
  and AND_11158(g22025,g5905,g19147);
  and AND_11159(g22026,g5913,g19147);
  and AND_11160(g22027,g5889,g19147);
  and AND_11161(g22028,g5893,g19147);
  and AND_11162(g22029,g5901,g19147);
  and AND_11163(g22030,g5909,g19147);
  and AND_11164(g22031,g5917,g19147);
  and AND_11165(g22032,g5921,g19147);
  and AND_11166(g22033,g5925,g19147);
  and AND_11167(g22034,g5929,g19147);
  and AND_11168(g22035,g5933,g19147);
  and AND_11169(g22036,g5937,g19147);
  and AND_11170(g22037,g5941,g19147);
  and AND_11171(g22038,g5945,g19147);
  and AND_11172(g22039,g5949,g19147);
  and AND_11173(g22040,g5953,g19147);
  and AND_11174(g22041,g5957,g19147);
  and AND_11175(g22042,g5961,g19147);
  and AND_11176(g22043,g5965,g19147);
  and AND_11177(g22044,g6058,g21611);
  and AND_11178(g22045,g6069,g21611);
  and AND_11179(g22046,g6073,g21611);
  and AND_11180(g22047,g6077,g21611);
  and AND_11181(g22048,g6052,g21611);
  and AND_11182(g22049,g6082,g21611);
  and AND_11183(g22050,g6088,g21611);
  and AND_11184(g22051,g6105,g21611);
  and AND_11185(g22052,g6113,g21611);
  and AND_11186(g22053,g6116,g21611);
  and AND_11187(g22054,g6120,g21611);
  and AND_11188(g22055,g6128,g21611);
  and AND_11189(g22056,g6133,g21611);
  and AND_11190(g22057,g15159,g21611);
  and AND_11191(g22058,g6098,g21611);
  and AND_11192(g22059,g6148,g21611);
  and AND_11193(g22060,g6151,g21611);
  and AND_11194(g22061,g6065,g21611);
  and AND_11195(g22062,g6093,g21611);
  and AND_11196(g22063,g6109,g21611);
  and AND_11197(g22064,g15162,g19210);
  and AND_11198(g22065,g6203,g19210);
  and AND_11199(g22066,g6209,g19210);
  and AND_11200(g22067,g6215,g19210);
  and AND_11201(g22068,g6219,g19210);
  and AND_11202(g22069,g6227,g19210);
  and AND_11203(g22070,g6243,g19210);
  and AND_11204(g22071,g6251,g19210);
  and AND_11205(g22072,g6259,g19210);
  and AND_11206(g22073,g6235,g19210);
  and AND_11207(g22074,g6239,g19210);
  and AND_11208(g22075,g6247,g19210);
  and AND_11209(g22076,g6255,g19210);
  and AND_11210(g22077,g6263,g19210);
  and AND_11211(g22078,g6267,g19210);
  and AND_11212(g22079,g6271,g19210);
  and AND_11213(g22080,g6275,g19210);
  and AND_11214(g22081,g6279,g19210);
  and AND_11215(g22082,g6283,g19210);
  and AND_11216(g22083,g6287,g19210);
  and AND_11217(g22084,g6291,g19210);
  and AND_11218(g22085,g6295,g19210);
  and AND_11219(g22086,g6299,g19210);
  and AND_11220(g22087,g6303,g19210);
  and AND_11221(g22088,g6307,g19210);
  and AND_11222(g22089,g6311,g19210);
  and AND_11223(g22090,g6404,g18833);
  and AND_11224(g22091,g6415,g18833);
  and AND_11225(g22092,g6419,g18833);
  and AND_11226(g22093,g6423,g18833);
  and AND_11227(g22094,g6398,g18833);
  and AND_11228(g22095,g6428,g18833);
  and AND_11229(g22096,g6434,g18833);
  and AND_11230(g22097,g6451,g18833);
  and AND_11231(g22098,g6459,g18833);
  and AND_11232(g22099,g6462,g18833);
  and AND_11233(g22100,g6466,g18833);
  and AND_11234(g22101,g6474,g18833);
  and AND_11235(g22102,g6479,g18833);
  and AND_11236(g22103,g15164,g18833);
  and AND_11237(g22104,g6444,g18833);
  and AND_11238(g22105,g6494,g18833);
  and AND_11239(g22106,g6497,g18833);
  and AND_11240(g22107,g6411,g18833);
  and AND_11241(g22108,g6439,g18833);
  and AND_11242(g22109,g6455,g18833);
  and AND_11243(g22110,g15167,g19277);
  and AND_11244(g22111,g6549,g19277);
  and AND_11245(g22112,g6555,g19277);
  and AND_11246(g22113,g6561,g19277);
  and AND_11247(g22114,g6565,g19277);
  and AND_11248(g22115,g6573,g19277);
  and AND_11249(g22116,g6589,g19277);
  and AND_11250(g22117,g6597,g19277);
  and AND_11251(g22118,g6605,g19277);
  and AND_11252(g22119,g6581,g19277);
  and AND_11253(g22120,g6585,g19277);
  and AND_11254(g22121,g6593,g19277);
  and AND_11255(g22122,g6601,g19277);
  and AND_11256(g22123,g6609,g19277);
  and AND_11257(g22124,g6613,g19277);
  and AND_11258(g22125,g6617,g19277);
  and AND_11259(g22126,g6621,g19277);
  and AND_11260(g22127,g6625,g19277);
  and AND_11261(g22128,g6629,g19277);
  and AND_11262(g22129,g6633,g19277);
  and AND_11263(g22130,g6637,g19277);
  and AND_11264(g22131,g6641,g19277);
  and AND_11265(g22132,g6645,g19277);
  and AND_11266(g22133,g6649,g19277);
  and AND_11267(g22134,g6653,g19277);
  and AND_11268(g22135,g6657,g19277);
  and AND_11269(g22142,g7957,g19140);
  and AND_11270(g22143,g19568,g10971);
  and AND_11271(g22145,g14555,g18832);
  and AND_11272(g22149,g14581,g18880);
  and AND_11273(g22157,g14608,g18892);
  and AND_11274(g22158,g13698,g19609);
  and AND_11275(g22160,g8005,g19795);
  and AND_11276(g22161,g13202,g19071);
  and AND_11277(g22165,g15594,g18903);
  and AND_11278(g22172,g8064,g19857);
  and AND_11279(g22191,g8119,g19875);
  and AND_11280(g22193,g19880,g20682);
  and AND_11281(g22208,g19906,g20739);
  and AND_11282(g22209,g19907,g20751);
  and AND_11283(g22216,g13660,g20000);
  and AND_11284(g22218,g19951,g20875);
  and AND_11285(g22219,g19953,g20887);
  and AND_11286(g22298,g19997,g21012);
  and AND_11287(g22299,g19999,g21024);
  and AND_11288(g22307,g20027,g21163);
  and AND_11289(g22308,g1135,g19738);
  and AND_11290(g22309,g1478,g19751);
  and AND_11291(g22310,g19662,g20235);
  and AND_11292(g22316,g2837,g20270);
  and AND_11293(g22329,g11940,g20329);
  and AND_11294(g22340,g19605,g13522);
  and AND_11295(g22342,g9354,g9285,g21287);
  and AND_11296(g22369,g9354,g7717,g20783);
  and AND_11297(g22384,g9354,g9285,g20784);
  and AND_11298(g22417,g7753,g9285,g21186);
  and AND_11299(g22432,g9354,g7717,g21187);
  and AND_11300(g22457,g7753,g7717,g21288);
  and AND_11301(g22472,g7753,g9285,g21289);
  and AND_11302(g22489,g12954,g19386);
  and AND_11303(g22498,g7753,g7717,g21334);
  and AND_11304(g22515,g12981,g19395);
  and AND_11305(g22518,g12982,g19398);
  and AND_11306(g22525,g13006,g19411);
  and AND_11307(g22534,g8766,g21389);
  and AND_11308(g22538,g14035,g20248);
  and AND_11309(g22588,g79,g20078);
  and AND_11310(g22589,g19267,g19451);
  and AND_11311(g22590,g19274,g19452);
  and AND_11312(g22622,g19336,g19469);
  and AND_11313(g22623,g19337,g19470);
  and AND_11314(g22624,g19344,g19471);
  and AND_11315(g22632,g19356,g19476);
  and AND_11316(g22633,g19359,g19479);
  and AND_11317(g22637,g19363,g19489);
  and AND_11318(g22665,g17174,g20905);
  and AND_11319(g22670,g20114,g9104);
  and AND_11320(g22680,g19530,g7781);
  and AND_11321(g22685,g11891,g20192);
  and AND_11322(g22686,g19335,g19577);
  and AND_11323(g22689,g18918,g9104);
  and AND_11324(g22710,g19358,g19600);
  and AND_11325(g22717,g9291,g20212);
  and AND_11326(g22720,g9253,g20619);
  and AND_11327(g22752,g15792,g19612);
  and AND_11328(g22760,g9360,g20237);
  and AND_11329(g22762,g9305,g20645);
  and AND_11330(g22831,g19441,g19629);
  and AND_11331(g22834,g102,g19630);
  and AND_11332(g22835,g15803,g19633);
  and AND_11333(g22843,g9429,g20272);
  and AND_11334(g22846,g9386,g20676);
  and AND_11335(g22848,g19449,g19649);
  and AND_11336(g22849,g1227,g19653);
  and AND_11337(g22851,g496,g19654);
  and AND_11338(g22859,g9456,g20734);
  and AND_11339(g22861,g19792,g19670);
  and AND_11340(g22862,g1570,g19673);
  and AND_11341(g22863,g9547,g20388);
  and AND_11342(g22871,g9523,g20871);
  and AND_11343(g22873,g19854,g19683);
  and AND_11344(g22876,g20136,g9104);
  and AND_11345(g22899,g19486,g19695);
  and AND_11346(g22900,g17137,g19697);
  and AND_11347(g22920,g19764,g19719);
  and AND_11348(g22937,g753,g20540);
  and AND_11349(g22938,g19782,g19739);
  and AND_11350(g22939,g9708,g21062);
  and AND_11351(g22942,g9104,g20219);
  and AND_11352(g22982,g19535,g19747);
  and AND_11353(g22990,g19555,g19760);
  and AND_11354(g22991,g645,g20248);
  and AND_11355(g22992,g1227,g19765);
  and AND_11356(g23006,g19575,g19776);
  and AND_11357(g23007,g681,g20248);
  and AND_11358(g23008,g1570,g19783);
  and AND_11359(g23009,g20196,g14219);
  and AND_11360(g23023,g650,g20248);
  and AND_11361(g23025,g16021,g19798);
  and AND_11362(g23050,g655,g20248);
  and AND_11363(g23056,g16052,g19860);
  and AND_11364(g23062,g718,g20248);
  and AND_11365(g23076,g19128,g9104);
  and AND_11366(g23083,g16076,g19878);
  and AND_11367(g23103,g10143,g20765);
  and AND_11368(g23104,g661,g20248);
  and AND_11369(g23121,g19128,g9104);
  and AND_11370(g23130,g728,g20248);
  and AND_11371(g23131,g13919,g19930);
  and AND_11372(g23148,g19128,g9104);
  and AND_11373(g23151,g18994,g7162);
  and AND_11374(g23165,g13954,g19964);
  and AND_11375(g23166,g13959,g19979);
  and AND_11376(g23187,g13989,g20010);
  and AND_11377(g23188,g13994,g20025);
  and AND_11378(g23201,g14027,g20040);
  and AND_11379(g23218,g20200,g16530);
  and AND_11380(g23220,g19417,g20067);
  and AND_11381(g23229,g18994,g4521);
  and AND_11382(g23254,g20056,g20110);
  and AND_11383(g23265,g20069,g20132);
  and AND_11384(g23280,g19417,g20146);
  and AND_11385(g23292,g19879,g16726);
  and AND_11386(g23293,g9104,g19200);
  and AND_11387(g23314,g9104,g19200);
  and AND_11388(g23348,g15570,g21393);
  and AND_11389(g23349,g13662,g20182);
  and AND_11390(g23372,g16448,g20194);
  and AND_11391(g23373,g13699,g20195);
  and AND_11392(g23381,g7239,g21413);
  and AND_11393(g23386,g20034,g20207);
  and AND_11394(g23387,g16506,g20211);
  and AND_11395(g23389,g9072,g19757);
  and AND_11396(g23392,g7247,g21430);
  and AND_11397(g23396,g20051,g20229);
  and AND_11398(g23397,g11154,g20239);
  and AND_11399(g23401,g7262,g21460);
  and AND_11400(g23404,g20063,g20247);
  and AND_11401(g23407,g9295,g20273);
  and AND_11402(g23412,g7297,g21510);
  and AND_11403(g23415,g20077,g20320);
  and AND_11404(g23416,g20082,g20321);
  and AND_11405(g23424,g7345,g21556);
  and AND_11406(g23436,g676,g20375);
  and AND_11407(g23439,g13771,g20452);
  and AND_11408(g23451,g13805,g20510);
  and AND_11409(g23471,g20148,g20523);
  and AND_11410(g23474,g13830,g20533);
  and AND_11411(g23475,g19070,g8971);
  and AND_11412(g23484,g20160,g20541);
  and AND_11413(g23497,g20169,g20569);
  and AND_11414(g23498,g20234,g12998);
  and AND_11415(g23513,g19430,g13007);
  and AND_11416(g23514,g20149,g11829);
  and AND_11417(g23531,g10760,g18930);
  and AND_11418(g23532,g19400,g11852);
  and AND_11419(g23533,g19436,g13015);
  and AND_11420(g23540,g16866,g20622);
  and AND_11421(g23551,g10793,g18948);
  and AND_11422(g23553,g19413,g11875);
  and AND_11423(g23554,g20390,g13024);
  and AND_11424(g23564,g16882,g20648);
  and AND_11425(g23572,g20230,g20656);
  and AND_11426(g23577,g19444,g13033);
  and AND_11427(g23581,g20183,g11900);
  and AND_11428(g23599,g19050,g9104);
  and AND_11429(g23606,g16927,g20679);
  and AND_11430(g23618,g19388,g11917);
  and AND_11431(g23619,g19453,g13045);
  and AND_11432(g23639,g19050,g9104);
  and AND_11433(g23646,g16959,g20737);
  and AND_11434(g23657,g19401,g11941);
  and AND_11435(g23658,g14687,g20852);
  and AND_11436(g23675,g19050,g9104);
  and AND_11437(g23682,g16970,g20874);
  and AND_11438(g23690,g14726,g20978);
  and AND_11439(g23691,g14731,g20993);
  and AND_11440(g23708,g19050,g9104);
  and AND_11441(g23724,g14767,g21123);
  and AND_11442(g23725,g14772,g21138);
  and AND_11443(g23742,g19128,g9104);
  and AND_11444(g23754,g14816,g21189);
  and AND_11445(g23755,g14821,g21204);
  and AND_11446(g23774,g14867,g21252);
  and AND_11447(g23775,g14872,g21267);
  and AND_11448(g23779,g1105,g19355);
  and AND_11449(g23799,g14911,g21279);
  and AND_11450(g23801,g1448,g19362);
  and AND_11451(g23802,g9104,g19050);
  and AND_11452(g23811,g4087,g19364);
  and AND_11453(g23828,g9104,g19128);
  and AND_11454(g23836,g4129,g19495);
  and AND_11455(g23837,g21160,g10804);
  and AND_11456(g23854,g4093,g19506);
  and AND_11457(g23855,g4112,g19455);
  and AND_11458(g23856,g4116,g19483);
  and AND_11459(g23857,g19626,g7908);
  and AND_11460(g23872,g19389,g4157);
  and AND_11461(g23873,g21222,g10815);
  and AND_11462(g23884,g4119,g19510);
  and AND_11463(g23885,g4132,g19513);
  and AND_11464(g23900,g1129,g19408);
  and AND_11465(g23901,g19606,g7963);
  and AND_11466(g23917,g1472,g19428);
  and AND_11467(g23919,g4122,g19546);
  and AND_11468(g23920,g4135,g19549);
  and AND_11469(g23921,g19379,g4146);
  and AND_11470(g23957,g4138,g19589);
  and AND_11471(g23958,g9104,g19200);
  and AND_11472(g23990,g19610,g10951);
  and AND_11473(g23991,g19209,g21428);
  and AND_11474(g23996,g19596,g10951);
  and AND_11475(g23998,g19631,g10971);
  and AND_11476(g24001,g19651,g10951);
  and AND_11477(g24002,g19613,g10971);
  and AND_11478(g24004,g37,g21225);
  and AND_11479(g24008,g7909,g19502);
  and AND_11480(g24009,g19671,g10971);
  and AND_11481(g24011,g7939,g19524);
  and AND_11482(g24012,g14496,g21561);
  and AND_11483(g24014,g7933,g19063);
  and AND_11484(g24015,g19540,g10951);
  and AND_11485(g24016,g14528,g21610);
  and AND_11486(g24139,g17619,g21653);
  and AND_11487(g24140,g17663,g21654);
  and AND_11488(g24141,g17657,g21656);
  and AND_11489(g24142,g17700,g21657);
  and AND_11490(g24143,g17694,g21659);
  and AND_11491(g24144,g17727,g21660);
  and AND_11492(g24186,g18102,g22722);
  and AND_11493(g24187,g305,g22722);
  and AND_11494(g24188,g316,g22722);
  and AND_11495(g24189,g324,g22722);
  and AND_11496(g24190,g329,g22722);
  and AND_11497(g24191,g319,g22722);
  and AND_11498(g24192,g311,g22722);
  and AND_11499(g24193,g336,g22722);
  and AND_11500(g24194,g106,g22722);
  and AND_11501(g24195,g74,g22722);
  and AND_11502(g24196,g333,g22722);
  and AND_11503(g24197,g347,g22722);
  and AND_11504(g24198,g351,g22722);
  and AND_11505(g24199,g355,g22722);
  and AND_11506(g24217,g18200,g22594);
  and AND_11507(g24218,g872,g22594);
  and AND_11508(g24219,g225,g22594);
  and AND_11509(g24220,g255,g22594);
  and AND_11510(g24221,g232,g22594);
  and AND_11511(g24222,g262,g22594);
  and AND_11512(g24223,g239,g22594);
  and AND_11513(g24224,g269,g22594);
  and AND_11514(g24225,g246,g22594);
  and AND_11515(g24226,g446,g22594);
  and AND_11516(g24227,g890,g22594);
  and AND_11517(g24228,g862,g22594);
  and AND_11518(g24229,g896,g22594);
  and AND_11519(g24230,g901,g22594);
  and AND_11520(g24283,g4411,g22550);
  and AND_11521(g24284,g4375,g22550);
  and AND_11522(g24285,g4388,g22550);
  and AND_11523(g24286,g4405,g22550);
  and AND_11524(g24287,g4401,g22550);
  and AND_11525(g24288,g4417,g22550);
  and AND_11526(g24289,g4427,g22550);
  and AND_11527(g24290,g4430,g22550);
  and AND_11528(g24291,g18660,g22550);
  and AND_11529(g24292,g4443,g22550);
  and AND_11530(g24293,g4438,g22550);
  and AND_11531(g24294,g4452,g22550);
  and AND_11532(g24295,g4434,g22550);
  and AND_11533(g24296,g4382,g22550);
  and AND_11534(g24297,g4455,g22550);
  and AND_11535(g24298,g4392,g22550);
  and AND_11536(g24299,g4456,g22550);
  and AND_11537(g24300,g15123,g22228);
  and AND_11538(g24301,g6961,g22228);
  and AND_11539(g24302,g15124,g22228);
  and AND_11540(g24303,g4369,g22228);
  and AND_11541(g24304,g12875,g22228);
  and AND_11542(g24305,g4477,g22228);
  and AND_11543(g24306,g4483,g22228);
  and AND_11544(g24307,g4486,g22228);
  and AND_11545(g24308,g4489,g22228);
  and AND_11546(g24309,g4480,g22228);
  and AND_11547(g24310,g4495,g22228);
  and AND_11548(g24311,g4498,g22228);
  and AND_11549(g24312,g4501,g22228);
  and AND_11550(g24313,g4504,g22228);
  and AND_11551(g24314,g4515,g22228);
  and AND_11552(g24315,g4521,g22228);
  and AND_11553(g24316,g4527,g22228);
  and AND_11554(g24317,g4534,g22228);
  and AND_11555(g24318,g4555,g22228);
  and AND_11556(g24319,g4561,g22228);
  and AND_11557(g24320,g6973,g22228);
  and AND_11558(g24321,g4558,g22228);
  and AND_11559(g24322,g4423,g22228);
  and AND_11560(g24323,g4546,g22228);
  and AND_11561(g24324,g4540,g22228);
  and AND_11562(g24325,g4543,g22228);
  and AND_11563(g24326,g4552,g22228);
  and AND_11564(g24327,g4549,g22228);
  and AND_11565(g24328,g4567,g22228);
  and AND_11566(g24329,g4462,g22228);
  and AND_11567(g24330,g18661,g22228);
  and AND_11568(g24331,g6977,g22228);
  and AND_11569(g24332,g4459,g22228);
  and AND_11570(g24333,g4512,g22228);
  and AND_11571(g24378,g3106,g22718);
  and AND_11572(g24387,g3457,g22761);
  and AND_11573(g24392,g3115,g23067);
  and AND_11574(g24393,g3808,g22844);
  and AND_11575(g24395,g4704,g22845);
  and AND_11576(g24399,g3133,g23067);
  and AND_11577(g24400,g3466,g23112);
  and AND_11578(g24402,g4749,g22857);
  and AND_11579(g24403,g4894,g22858);
  and AND_11580(g24406,g13623,g22860);
  and AND_11581(g24408,g23989,g18946);
  and AND_11582(g24409,g3484,g23112);
  and AND_11583(g24410,g3817,g23139);
  and AND_11584(g24411,g4584,g22161);
  and AND_11585(g24415,g4760,g22869);
  and AND_11586(g24416,g4939,g22870);
  and AND_11587(g24420,g23997,g18980);
  and AND_11588(g24421,g3835,g23139);
  and AND_11589(g24422,g4771,g22896);
  and AND_11590(g24423,g4950,g22897);
  and AND_11591(g24427,g4961,g22919);
  and AND_11592(g24436,g3125,g23067);
  and AND_11593(g24450,g3129,g23067);
  and AND_11594(g24451,g3476,g23112);
  and AND_11595(g24464,g3480,g23112);
  and AND_11596(g24465,g3827,g23139);
  and AND_11597(g24467,g13761,g23047);
  and AND_11598(g24475,g3831,g23139);
  and AND_11599(g24476,g18879,g22330);
  and AND_11600(g24482,g6875,g23055);
  and AND_11601(g24484,g16288,g23208);
  and AND_11602(g24485,g10710,g22319);
  and AND_11603(g24488,g6905,g23082);
  and AND_11604(g24491,g10727,g22332);
  and AND_11605(g24495,g6928,g23127);
  and AND_11606(g24498,g14036,g23850);
  and AND_11607(g24499,g22217,g19394);
  and AND_11608(g24501,g14000,g23182);
  and AND_11609(g24502,g23428,g13223);
  and AND_11610(g24503,g22225,g19409);
  and AND_11611(g24504,g22226,g19410);
  and AND_11612(g24507,g22304,g19429);
  and AND_11613(g24523,g22318,g19468);
  and AND_11614(g24532,g22331,g19478);
  and AND_11615(g24536,g19516,g22635);
  and AND_11616(g24537,g22626,g10851);
  and AND_11617(g24541,g22626,g10851);
  and AND_11618(g24545,g3333,g23285);
  and AND_11619(g24546,g22447,g19523);
  and AND_11620(g24549,g23162,g20887);
  and AND_11621(g24550,g3684,g23308);
  and AND_11622(g24551,g17148,g23331);
  and AND_11623(g24552,g22487,g19538);
  and AND_11624(g24553,g22983,g19539);
  and AND_11625(g24554,g22490,g19541);
  and AND_11626(g24555,g23184,g21024);
  and AND_11627(g24556,g4035,g23341);
  and AND_11628(g24558,g22516,g19566);
  and AND_11629(g24559,g22993,g19567);
  and AND_11630(g24564,g23198,g21163);
  and AND_11631(g24569,g5115,g23382);
  and AND_11632(g24572,g5462,g23393);
  and AND_11633(g24573,g17198,g23716);
  and AND_11634(g24581,g5124,g23590);
  and AND_11635(g24582,g5808,g23402);
  and AND_11636(g24588,g5142,g23590);
  and AND_11637(g24589,g5471,g23630);
  and AND_11638(g24590,g6154,g23413);
  and AND_11639(g24600,g22591,g19652);
  and AND_11640(g24602,g16507,g22854);
  and AND_11641(g24606,g5489,g23630);
  and AND_11642(g24607,g5817,g23666);
  and AND_11643(g24608,g6500,g23425);
  and AND_11644(g24618,g22625,g19672);
  and AND_11645(g24622,g19856,g22866);
  and AND_11646(g24624,g16524,g22867);
  and AND_11647(g24627,g22763,g19679);
  and AND_11648(g24628,g5835,g23666);
  and AND_11649(g24629,g6163,g23699);
  and AND_11650(g24630,g23255,g14149);
  and AND_11651(g24634,g22634,g19685);
  and AND_11652(g24635,g19874,g22883);
  and AND_11653(g24637,g16586,g22884);
  and AND_11654(g24638,g22763,g19690);
  and AND_11655(g24639,g6181,g23699);
  and AND_11656(g24640,g6509,g23733);
  and AND_11657(g24642,g8290,g22898);
  and AND_11658(g24643,g22636,g19696);
  and AND_11659(g24644,g11714,g22903);
  and AND_11660(g24645,g22639,g19709);
  and AND_11661(g24646,g22640,g19711);
  and AND_11662(g24647,g19903,g22907);
  and AND_11663(g24649,g6527,g23733);
  and AND_11664(g24650,g22641,g19718);
  and AND_11665(g24651,g2741,g23472);
  and AND_11666(g24654,g11735,g22922);
  and AND_11667(g24656,g11736,g22926);
  and AND_11668(g24657,g22644,g19730);
  and AND_11669(g24658,g22645,g19732);
  and AND_11670(g24659,g5134,g23590);
  and AND_11671(g24660,g22648,g19737);
  and AND_11672(g24663,g16621,g22974);
  and AND_11673(g24664,g22652,g19741);
  and AND_11674(g24666,g11753,g22975);
  and AND_11675(g24668,g11754,g22979);
  and AND_11676(g24669,g22653,g19742);
  and AND_11677(g24670,g5138,g23590);
  and AND_11678(g24671,g5481,g23630);
  and AND_11679(g24672,g19534,g22981);
  and AND_11680(g24673,g22659,g19748);
  and AND_11681(g24674,g446,g23496);
  and AND_11682(g24675,g17568,g22342);
  and AND_11683(g24676,g2748,g23782);
  and AND_11684(g24679,g13289,g22985);
  and AND_11685(g24680,g16422,g22986);
  and AND_11686(g24681,g16653,g22988);
  and AND_11687(g24682,g22662,g19754);
  and AND_11688(g24684,g11769,g22989);
  and AND_11689(g24686,g5485,g23630);
  and AND_11690(g24687,g5827,g23666);
  and AND_11691(g24688,g22681,g22663);
  and AND_11692(g24698,g22664,g19761);
  and AND_11693(g24700,g645,g23512);
  and AND_11694(g24702,g17464,g22342);
  and AND_11695(g24703,g17592,g22369);
  and AND_11696(g24704,g17593,g22384);
  and AND_11697(g24706,g15910,g22996);
  and AND_11698(g24707,g13295,g22997);
  and AND_11699(g24708,g16474,g22998);
  and AND_11700(g24709,g16690,g23000);
  and AND_11701(g24710,g22679,g19771);
  and AND_11702(g24712,g19592,g23001);
  and AND_11703(g24713,g5831,g23666);
  and AND_11704(g24714,g6173,g23699);
  and AND_11705(g24716,g15935,g23004);
  and AND_11706(g24717,g22684,g19777);
  and AND_11707(g24719,g681,g23530);
  and AND_11708(g24721,g17488,g22369);
  and AND_11709(g24722,g17618,g22417);
  and AND_11710(g24723,g17490,g22384);
  and AND_11711(g24724,g17624,g22432);
  and AND_11712(g24725,g19587,g23012);
  and AND_11713(g24726,g15965,g23015);
  and AND_11714(g24727,g13300,g23016);
  and AND_11715(g24728,g16513,g23017);
  and AND_11716(g24729,g22719,g23018);
  and AND_11717(g24730,g6177,g23699);
  and AND_11718(g24731,g6519,g23733);
  and AND_11719(g24743,g22708,g19789);
  and AND_11720(g24745,g650,g23550);
  and AND_11721(g24747,g17510,g22417);
  and AND_11722(g24748,g17656,g22457);
  and AND_11723(g24749,g17511,g22432);
  and AND_11724(g24750,g17662,g22472);
  and AND_11725(g24754,g19604,g23027);
  and AND_11726(g24755,g16022,g23030);
  and AND_11727(g24757,g7004,g23563);
  and AND_11728(g24758,g6523,g23733);
  and AND_11729(g24761,g22751,g19852);
  and AND_11730(g24762,g655,g23573);
  and AND_11731(g24763,g17569,g22457);
  and AND_11732(g24764,g17570,g22472);
  and AND_11733(g24765,g17699,g22498);
  and AND_11734(g24769,g19619,g23058);
  and AND_11735(g24771,g7028,g23605);
  and AND_11736(g24772,g16287,g23061);
  and AND_11737(g24773,g22832,g19872);
  and AND_11738(g24774,g718,g23614);
  and AND_11739(g24775,g17594,g22498);
  and AND_11740(g24777,g11345,g23066);
  and AND_11741(g24785,g7051,g23645);
  and AND_11742(g24786,g661,g23654);
  and AND_11743(g24788,g11384,g23111);
  and AND_11744(g24790,g7074,g23681);
  and AND_11745(g24794,g11414,g23138);
  and AND_11746(g24796,g7097,g23714);
  and AND_11747(g24797,g22872,g19960);
  and AND_11748(g24803,g22901,g20005);
  and AND_11749(g24812,g19662,g22192);
  and AND_11750(g24817,g22929,g7235);
  and AND_11751(g24820,g13944,g23978);
  and AND_11752(I24003,g8097,g8334,g3045);
  and AND_11753(g24822,g3010,g23534,I24003);
  and AND_11754(g24835,g8720,g23233);
  and AND_11755(I24015,g8334,g7975,g3045);
  and AND_11756(g24843,g3010,g23211,I24015);
  and AND_11757(I24018,g8155,g8390,g3396);
  and AND_11758(g24846,g3361,g23555,I24018);
  and AND_11759(g24849,g4165,g22227);
  and AND_11760(I24027,g3029,g3034,g8426);
  and AND_11761(g24855,g3050,g23534,I24027);
  and AND_11762(I24030,g8390,g8016,g3396);
  and AND_11763(g24858,g3361,g23223,I24030);
  and AND_11764(I24033,g8219,g8443,g3747);
  and AND_11765(g24861,g3712,g23582,I24033);
  and AND_11766(g24864,g11201,g22305);
  and AND_11767(g24865,g11323,g23253);
  and AND_11768(g24872,g23088,g9104);
  and AND_11769(I24048,g3034,g3040,g8426);
  and AND_11770(g24881,g3050,g23211,I24048);
  and AND_11771(I24051,g3380,g3385,g8492);
  and AND_11772(g24884,g3401,g23555,I24051);
  and AND_11773(I24054,g8443,g8075,g3747);
  and AND_11774(g24887,g3712,g23239,I24054);
  and AND_11775(g24892,g11559,g23264);
  and AND_11776(I24064,g3385,g3391,g8492);
  and AND_11777(g24897,g3401,g23223,I24064);
  and AND_11778(I24067,g3731,g3736,g8553);
  and AND_11779(g24900,g3752,g23582,I24067);
  and AND_11780(g24903,g128,g23889);
  and AND_11781(g24904,g11761,g23279);
  and AND_11782(I24075,g3736,g3742,g8553);
  and AND_11783(g24908,g3752,g23239,I24075);
  and AND_11784(g24912,g23687,g20682);
  and AND_11785(g24913,g4821,g23908);
  and AND_11786(g24914,g8721,g23301);
  and AND_11787(g24915,g23087,g20158);
  and AND_11788(g24921,g23721,g20739);
  and AND_11789(g24922,g4831,g23931);
  and AND_11790(g24923,g23129,g20167);
  and AND_11791(g24929,g23751,g20875);
  and AND_11792(g24930,g4826,g23948);
  and AND_11793(g24931,g23153,g20178);
  and AND_11794(g24939,g23771,g21012);
  and AND_11795(g24940,g5011,g23971);
  and AND_11796(g24941,g23171,g20190);
  and AND_11797(g24945,g23183,g20197);
  and AND_11798(g24949,g23796,g20751);
  and AND_11799(g24961,g23193,g20209);
  and AND_11800(g24962,g23194,g20210);
  and AND_11801(g24967,g23197,g20213);
  and AND_11802(g24977,g23209,g20232);
  and AND_11803(g24983,g23217,g20238);
  and AND_11804(g24984,g22929,g12818);
  and AND_11805(g24997,g22929,g10419);
  and AND_11806(g24998,g17412,g23408);
  and AND_11807(g25012,g20644,g23419);
  and AND_11808(g25014,g17474,g23420);
  and AND_11809(g25026,g22929,g10503);
  and AND_11810(g25030,g23251,g20432);
  and AND_11811(g25031,g20675,g23432);
  and AND_11812(g25033,g17500,g23433);
  and AND_11813(g25040,g12738,g23443);
  and AND_11814(g25041,g23261,g20494);
  and AND_11815(g25042,g23262,g20496);
  and AND_11816(g25043,g20733,g23447);
  and AND_11817(g25045,g17525,g23448);
  and AND_11818(g25050,g13056,g22312);
  and AND_11819(g25054,g12778,g23452);
  and AND_11820(g25056,g12779,g23456);
  and AND_11821(g25057,g23275,g20511);
  and AND_11822(g25058,g23276,g20513);
  and AND_11823(g25059,g20870,g23460);
  and AND_11824(g25061,g17586,g23461);
  and AND_11825(g25063,g13078,g22325);
  and AND_11826(g25067,g4722,g22885);
  and AND_11827(g25068,g17574,g23477);
  and AND_11828(g25069,g23296,g20535);
  and AND_11829(g25071,g12804,g23478);
  and AND_11830(g25076,g12805,g23479);
  and AND_11831(g25077,g23297,g20536);
  and AND_11832(g25078,g23298,g20538);
  and AND_11833(g25079,g21011,g23483);
  and AND_11834(g25084,g4737,g22885);
  and AND_11835(g25085,g4912,g22908);
  and AND_11836(g25086,g13941,g23488);
  and AND_11837(g25087,g17307,g23489);
  and AND_11838(g25088,g17601,g23491);
  and AND_11839(g25089,g23317,g20553);
  and AND_11840(g25091,g12830,g23492);
  and AND_11841(g25093,g12831,g23493);
  and AND_11842(g25094,g23318,g20554);
  and AND_11843(g25095,g23319,g20556);
  and AND_11844(g25096,g23778,g20560);
  and AND_11845(g25102,g4727,g22885);
  and AND_11846(g25103,g4927,g22908);
  and AND_11847(g25104,g16800,g23504);
  and AND_11848(g25105,g13973,g23505);
  and AND_11849(g25106,g17391,g23506);
  and AND_11850(g25107,g17643,g23508);
  and AND_11851(g25108,g23345,g20576);
  and AND_11852(g25110,g10427,g23509);
  and AND_11853(g25112,g10428,g23510);
  and AND_11854(g25113,g23346,g20577);
  and AND_11855(g25122,g23374,g20592);
  and AND_11856(g25123,g4732,g22885);
  and AND_11857(g25124,g4917,g22908);
  and AND_11858(g25125,g20187,g23520);
  and AND_11859(g25126,g16839,g23523);
  and AND_11860(g25127,g13997,g23524);
  and AND_11861(g25128,g17418,g23525);
  and AND_11862(g25129,g17682,g23527);
  and AND_11863(g25130,g23358,g20600);
  and AND_11864(g25132,g10497,g23528);
  and AND_11865(g25142,g4717,g22885);
  and AND_11866(g25143,g4922,g22908);
  and AND_11867(g25147,g20202,g23542);
  and AND_11868(g25148,g16867,g23545);
  and AND_11869(g25149,g14030,g23546);
  and AND_11870(g25150,g17480,g23547);
  and AND_11871(g25151,g17719,g23549);
  and AND_11872(g25152,g23383,g20626);
  and AND_11873(g25159,g4907,g22908);
  and AND_11874(g25163,g20217,g23566);
  and AND_11875(g25164,g16883,g23569);
  and AND_11876(g25165,g14062,g23570);
  and AND_11877(g25166,g17506,g23571);
  and AND_11878(g25173,g12234,g23589);
  and AND_11879(g25178,g20241,g23608);
  and AND_11880(g25179,g16928,g23611);
  and AND_11881(g25181,g23405,g20696);
  and AND_11882(g25187,g12296,g23629);
  and AND_11883(g25192,g20276,g23648);
  and AND_11884(g25201,g12346,g23665);
  and AND_11885(g25207,g22513,g10621);
  and AND_11886(g25217,g12418,g23698);
  and AND_11887(g25223,g22523,g10652);
  and AND_11888(g25229,g7636,g22654);
  and AND_11889(g25238,g12466,g23732);
  and AND_11890(g25285,g22152,g13061);
  and AND_11891(I24482,g9364,g9607,g5057);
  and AND_11892(g25290,g5022,g22173,I24482);
  and AND_11893(g25323,g6888,g22359);
  and AND_11894(I24505,g9607,g9229,g5057);
  and AND_11895(g25328,g5022,g23764,I24505);
  and AND_11896(I24508,g9434,g9672,g5401);
  and AND_11897(g25331,g5366,g22194,I24508);
  and AND_11898(g25357,g23810,g23786);
  and AND_11899(g25366,g7733,g22406);
  and AND_11900(g25367,g6946,g22407);
  and AND_11901(g25368,g6946,g22408);
  and AND_11902(I24524,g5041,g5046,g9716);
  and AND_11903(g25371,g5062,g22173,I24524);
  and AND_11904(I24527,g9672,g9264,g5401);
  and AND_11905(g25374,g5366,g23789,I24527);
  and AND_11906(I24530,g9501,g9733,g5747);
  and AND_11907(g25377,g5712,g22210,I24530);
  and AND_11908(g25408,g22682,g9772);
  and AND_11909(I24546,g5046,g5052,g9716);
  and AND_11910(g25411,g5062,g23764,I24546);
  and AND_11911(I24549,g5385,g5390,g9792);
  and AND_11912(g25414,g5406,g22194,I24549);
  and AND_11913(I24552,g9733,g9316,g5747);
  and AND_11914(g25417,g5712,g23816,I24552);
  and AND_11915(I24555,g9559,g9809,g6093);
  and AND_11916(g25420,g6058,g22220,I24555);
  and AND_11917(g25448,g11202,g22680);
  and AND_11918(g25449,g6946,g22496);
  and AND_11919(g25450,g6888,g22497);
  and AND_11920(I24576,g5390,g5396,g9792);
  and AND_11921(g25453,g5406,g23789,I24576);
  and AND_11922(I24579,g5731,g5736,g9875);
  and AND_11923(g25456,g5752,g22210,I24579);
  and AND_11924(I24582,g9809,g9397,g6093);
  and AND_11925(g25459,g6058,g23844,I24582);
  and AND_11926(I24585,g9621,g9892,g6439);
  and AND_11927(g25462,g6404,g22300,I24585);
  and AND_11928(g25466,g23574,g21346);
  and AND_11929(g25479,g22646,g9917);
  and AND_11930(I24597,g5736,g5742,g9875);
  and AND_11931(g25482,g5752,g23816,I24597);
  and AND_11932(I24600,g6077,g6082,g9946);
  and AND_11933(g25485,g6098,g22220,I24600);
  and AND_11934(I24603,g9892,g9467,g6439);
  and AND_11935(g25488,g6404,g23865,I24603);
  and AND_11936(g25491,g23615,g21355);
  and AND_11937(g25502,g6946,g22527);
  and AND_11938(g25503,g6888,g22529);
  and AND_11939(I24616,g6082,g6088,g9946);
  and AND_11940(g25507,g6098,g23844,I24616);
  and AND_11941(I24619,g6423,g6428,g10014);
  and AND_11942(g25510,g6444,g22300,I24619);
  and AND_11943(I24625,g6428,g6434,g10014);
  and AND_11944(g25518,g6444,g23865,I24625);
  and AND_11945(g25522,g6888,g22544);
  and AND_11946(g25526,g23720,g21400);
  and AND_11947(g25530,g23750,g21414);
  and AND_11948(g25536,g23770,g21431);
  and AND_11949(g25543,g23795,g21461);
  and AND_11950(g25551,g23822,g21511);
  and AND_11951(g25559,g13004,g22649);
  and AND_11952(g25565,g13013,g22660);
  and AND_11953(I24674,g19919,g24019,g24020,g24021);
  and AND_11954(I24675,g24022,g24023,g24024,g24025);
  and AND_11955(g25567,I24674,I24675);
  and AND_11956(I24679,g19968,g24026,g24027,g24028);
  and AND_11957(I24680,g24029,g24030,g24031,g24032);
  and AND_11958(g25568,I24679,I24680);
  and AND_11959(I24684,g20014,g24033,g24034,g24035);
  and AND_11960(I24685,g24036,g24037,g24038,g24039);
  and AND_11961(g25569,I24684,I24685);
  and AND_11962(I24689,g20841,g24040,g24041,g24042);
  and AND_11963(I24690,g24043,g24044,g24045,g24046);
  and AND_11964(g25570,I24689,I24690);
  and AND_11965(I24694,g20982,g24047,g24048,g24049);
  and AND_11966(I24695,g24050,g24051,g24052,g24053);
  and AND_11967(g25571,I24694,I24695);
  and AND_11968(I24699,g21127,g24054,g24055,g24056);
  and AND_11969(I24700,g24057,g24058,g24059,g24060);
  and AND_11970(g25572,I24699,I24700);
  and AND_11971(I24704,g21193,g24061,g24062,g24063);
  and AND_11972(I24705,g24064,g24065,g24066,g24067);
  and AND_11973(g25573,I24704,I24705);
  and AND_11974(I24709,g21256,g24068,g24069,g24070);
  and AND_11975(I24710,g24071,g24072,g24073,g24074);
  and AND_11976(g25574,I24709,I24710);
  and AND_11977(g25578,g19402,g24146);
  and AND_11978(g25579,g19422,g24147);
  and AND_11979(g25580,g19268,g24149);
  and AND_11980(g25581,g19338,g24150);
  and AND_11981(g25765,g24989,g24973);
  and AND_11982(g25768,g2912,g24560);
  and AND_11983(g25772,g24944,g24934);
  and AND_11984(g25775,g2922,g24568);
  and AND_11985(g25780,g25532,g25527);
  and AND_11986(g25782,g2936,g24571);
  and AND_11987(g25787,g24792,g20887);
  and AND_11988(g25788,g8010,g24579);
  and AND_11989(g25801,g8097,g24585);
  and AND_11990(g25802,g8106,g24586);
  and AND_11991(g25803,g24798,g21024);
  and AND_11992(g25804,g8069,g24587);
  and AND_11993(g25814,g24760,g13323);
  and AND_11994(g25815,g8155,g24603);
  and AND_11995(g25816,g8164,g24604);
  and AND_11996(g25817,g24807,g21163);
  and AND_11997(g25818,g8124,g24605);
  and AND_11998(g25831,g3151,g24623);
  and AND_11999(g25832,g8219,g24625);
  and AND_12000(g25833,g8228,g24626);
  and AND_12001(g25848,g25539,g18977);
  and AND_12002(g25850,g3502,g24636);
  and AND_12003(g25852,g4593,g24411);
  and AND_12004(g25865,g25545,g18991);
  and AND_12005(g25866,g3853,g24648);
  and AND_12006(g25870,g24840,g16182);
  and AND_12007(g25871,g8334,g24804);
  and AND_12008(g25872,g3119,g24655);
  and AND_12009(g25873,g24854,g16197);
  and AND_12010(g25874,g11118,g24665);
  and AND_12011(g25875,g8390,g24809);
  and AND_12012(g25876,g3470,g24667);
  and AND_12013(g25879,g11135,g24683);
  and AND_12014(g25880,g8443,g24814);
  and AND_12015(g25881,g3821,g24685);
  and AND_12016(g25883,g13728,g24699);
  and AND_12017(g25884,g11153,g24711);
  and AND_12018(g25900,g24390,g19368);
  and AND_12019(g25901,g24853,g16290);
  and AND_12020(g25902,g24398,g19373);
  and AND_12021(g25904,g14001,g24791);
  and AND_12022(g25905,g24879,g16311);
  and AND_12023(g25907,g24799,g22519);
  and AND_12024(g25908,g24782,g22520);
  and AND_12025(g25909,g8745,g24875);
  and AND_12026(g25915,g24926,g9602);
  and AND_12027(g25916,g24432,g19434);
  and AND_12028(g25921,g24936,g9664);
  and AND_12029(g25922,g24959,g20065);
  and AND_12030(g25923,g24443,g19443);
  and AND_12031(g25924,g24976,g16846);
  and AND_12032(g25925,g24990,g23234);
  and AND_12033(g25926,g25005,g24839);
  and AND_12034(g25927,g25004,g20375);
  and AND_12035(g25928,g25022,g23436);
  and AND_12036(g25931,g24574,g19477);
  and AND_12037(g25938,g8997,g24953);
  and AND_12038(g25939,g24583,g19490);
  and AND_12039(g25946,g24496,g19537);
  and AND_12040(g25949,g24701,g19559);
  and AND_12041(g25951,g24500,g19565);
  and AND_12042(g25955,g24720,g19580);
  and AND_12043(g25957,g17190,g24960);
  and AND_12044(g25959,g1648,g24963);
  and AND_12045(g25961,g25199,g20682);
  and AND_12046(g25962,g9258,g24971);
  and AND_12047(g25963,g1657,g24978);
  and AND_12048(g25964,g1783,g24979);
  and AND_12049(g25965,g2208,g24980);
  and AND_12050(g25966,g9364,g24985);
  and AND_12051(g25967,g9373,g24986);
  and AND_12052(g25968,g25215,g20739);
  and AND_12053(g25969,g9310,g24987);
  and AND_12054(g25970,g1792,g24991);
  and AND_12055(g25971,g1917,g24992);
  and AND_12056(g25972,g2217,g24993);
  and AND_12057(g25973,g2342,g24994);
  and AND_12058(g25975,g9434,g24999);
  and AND_12059(g25976,g9443,g25000);
  and AND_12060(g25977,g25236,g20875);
  and AND_12061(g25978,g9391,g25001);
  and AND_12062(g25979,g24517,g19650);
  and AND_12063(g25980,g1926,g25006);
  and AND_12064(g25981,g2051,g25007);
  and AND_12065(g25982,g2351,g25008);
  and AND_12066(g25983,g2476,g25009);
  and AND_12067(g25986,g5160,g25013);
  and AND_12068(g25987,g9501,g25015);
  and AND_12069(g25988,g9510,g25016);
  and AND_12070(g25989,g25258,g21012);
  and AND_12071(g25990,g9461,g25017);
  and AND_12072(g25991,g2060,g25023);
  and AND_12073(g25992,g2485,g25024);
  and AND_12074(g25993,g2610,g25025);
  and AND_12075(g26019,g5507,g25032);
  and AND_12076(g26020,g9559,g25034);
  and AND_12077(g26021,g9568,g25035);
  and AND_12078(g26022,g25271,g20751);
  and AND_12079(g26023,g9528,g25036);
  and AND_12080(g26024,g2619,g25039);
  and AND_12081(g26048,g5853,g25044);
  and AND_12082(g26049,g9621,g25046);
  and AND_12083(g26050,g9630,g25047);
  and AND_12084(g26051,g24896,g14169);
  and AND_12085(g26077,g9607,g25233);
  and AND_12086(g26078,g5128,g25055);
  and AND_12087(g26079,g6199,g25060);
  and AND_12088(g26084,g24926,g9602);
  and AND_12089(g26085,g11906,g25070);
  and AND_12090(g26086,g9672,g25255);
  and AND_12091(g26087,g5475,g25072);
  and AND_12092(g26088,g6545,g25080);
  and AND_12093(g26090,g1624,g25081);
  and AND_12094(g26091,g1691,g25082);
  and AND_12095(g26092,g9766,g25083);
  and AND_12096(g26094,g24936,g9664);
  and AND_12097(g26095,g11923,g25090);
  and AND_12098(g26096,g9733,g25268);
  and AND_12099(g26097,g5821,g25092);
  and AND_12100(g26100,g1677,g25097);
  and AND_12101(g26101,g1760,g25098);
  and AND_12102(g26102,g1825,g25099);
  and AND_12103(g26103,g2185,g25100);
  and AND_12104(g26104,g2250,g25101);
  and AND_12105(g26119,g11944,g25109);
  and AND_12106(g26120,g9809,g25293);
  and AND_12107(g26121,g6167,g25111);
  and AND_12108(g26122,g24557,g19762);
  and AND_12109(g26123,g1696,g25382);
  and AND_12110(g26124,g1811,g25116);
  and AND_12111(g26125,g1894,g25117);
  and AND_12112(g26126,g1959,g25118);
  and AND_12113(g26127,g2236,g25119);
  and AND_12114(g26128,g2319,g25120);
  and AND_12115(g26129,g2384,g25121);
  and AND_12116(g26130,g24890,g19772);
  and AND_12117(g26145,g11962,g25131);
  and AND_12118(g26146,g9892,g25334);
  and AND_12119(g26147,g6513,g25133);
  and AND_12120(g26148,g25357,g11724,g11709,g11686);
  and AND_12121(g26153,g24565,g19780);
  and AND_12122(g26154,g1830,g25426);
  and AND_12123(g26155,g1945,g25134);
  and AND_12124(g26156,g2028,g25135);
  and AND_12125(g26157,g2093,g25136);
  and AND_12126(g26158,g2255,g25432);
  and AND_12127(g26159,g2370,g25137);
  and AND_12128(g26160,g2453,g25138);
  and AND_12129(g26161,g2518,g25139);
  and AND_12130(g26165,g11980,g25153);
  and AND_12131(g26166,g25357,g11724,g11709,g7558);
  and AND_12132(g26171,g25357,g6856,g11709,g11686);
  and AND_12133(g26176,g1964,g25467);
  and AND_12134(g26177,g2079,g25154);
  and AND_12135(g26178,g2389,g25473);
  and AND_12136(g26179,g2504,g25155);
  and AND_12137(g26180,g2587,g25156);
  and AND_12138(g26181,g2652,g25157);
  and AND_12139(g26182,g9978,g25317);
  and AND_12140(g26186,g24580,g23031);
  and AND_12141(g26190,g25357,g11724,g7586,g11686);
  and AND_12142(g26195,g25357,g6856,g11709,g7558);
  and AND_12143(g26200,g24688,g10678,g10658,g10627);
  and AND_12144(g26203,g1632,g25337);
  and AND_12145(g26204,g1720,g25275);
  and AND_12146(g26205,g2098,g25492);
  and AND_12147(g26206,g2523,g25495);
  and AND_12148(g26207,g2638,g25170);
  and AND_12149(g26213,g25357,g11724,g7586,g7558);
  and AND_12150(g26218,g25357,g6856,g7586,g11686);
  and AND_12151(g26223,g24688,g10678,g10658,g8757);
  and AND_12152(g26226,g24688,g8812,g10658,g10627);
  and AND_12153(g26229,g1724,g25275);
  and AND_12154(g26230,g1768,g25385);
  and AND_12155(g26231,g1854,g25300);
  and AND_12156(g26232,g2193,g25396);
  and AND_12157(g26233,g2279,g25309);
  and AND_12158(g26234,g2657,g25514);
  and AND_12159(g26236,g25357,g6856,g7586,g7558);
  and AND_12160(g26241,g24688,g10678,g8778,g10627);
  and AND_12161(g26244,g24688,g8812,g10658,g8757);
  and AND_12162(g26249,g1858,g25300);
  and AND_12163(g26250,g1902,g25429);
  and AND_12164(g26251,g1988,g25341);
  and AND_12165(g26252,g2283,g25309);
  and AND_12166(g26253,g2327,g25435);
  and AND_12167(g26254,g2413,g25349);
  and AND_12168(g26257,g4253,g25197);
  and AND_12169(g26258,g12875,g25231);
  and AND_12170(g26259,g24430,g25232);
  and AND_12171(g26261,g24688,g10678,g8778,g8757);
  and AND_12172(g26264,g24688,g8812,g8778,g10627);
  and AND_12173(g26270,g1700,g25275);
  and AND_12174(g26271,g1992,g25341);
  and AND_12175(g26272,g2036,g25470);
  and AND_12176(g26273,g2122,g25389);
  and AND_12177(g26274,g2130,g25210);
  and AND_12178(g26275,g2417,g25349);
  and AND_12179(g26276,g2461,g25476);
  and AND_12180(g26277,g2547,g25400);
  and AND_12181(g26279,g4249,g25213);
  and AND_12182(g26280,g13051,g25248);
  and AND_12183(g26281,g24688,g8812,g8778,g8757);
  and AND_12184(g26285,g1834,g25300);
  and AND_12185(g26286,g2126,g25389);
  and AND_12186(g26287,g2138,g25225);
  and AND_12187(g26288,g2259,g25309);
  and AND_12188(g26289,g2551,g25400);
  and AND_12189(g26290,g2595,g25498);
  and AND_12190(g26291,g2681,g25439);
  and AND_12191(g26292,g2689,g25228);
  and AND_12192(g26294,g4245,g25230);
  and AND_12193(g26295,g13070,g25266);
  and AND_12194(g26300,g1968,g25341);
  and AND_12195(g26301,g2145,g25244);
  and AND_12196(g26302,g2393,g25349);
  and AND_12197(g26303,g2685,g25439);
  and AND_12198(g26304,g2697,g25246);
  and AND_12199(g26306,g13087,g25286);
  and AND_12200(g26307,g13070,g25288);
  and AND_12201(g26308,g6961,g25289);
  and AND_12202(g26310,g2102,g25389);
  and AND_12203(g26311,g2527,g25400);
  and AND_12204(g26312,g2704,g25264);
  and AND_12205(g26313,g12645,g25326);
  and AND_12206(g26323,g10262,g25273);
  and AND_12207(g26324,g2661,g25439);
  and AND_12208(g26325,g12644,g25370);
  and AND_12209(g26336,g10307,g25480);
  and AND_12210(g26339,g225,g24836);
  and AND_12211(g26341,g24746,g20105);
  and AND_12212(g26345,g13051,g25505);
  and AND_12213(g26347,g262,g24850);
  and AND_12214(g26350,g13087,g25517);
  and AND_12215(g26351,g239,g24869);
  and AND_12216(g26356,g15581,g25523);
  and AND_12217(g26357,g22547,g25525);
  and AND_12218(g26358,g19522,g25528);
  and AND_12219(g26360,g10589,g25533);
  and AND_12220(g26362,g19557,g25538);
  and AND_12221(g26378,g19576,g25544);
  and AND_12222(g26379,g19904,g25546);
  and AND_12223(g26380,g19572,g25547);
  and AND_12224(g26381,g4456,g25548);
  and AND_12225(g26387,g24813,g20231);
  and AND_12226(g26388,g19595,g25552);
  and AND_12227(g26389,g19949,g25553);
  and AND_12228(g26390,g4423,g25554);
  and AND_12229(g26391,g19593,g25555);
  and AND_12230(g26393,g19467,g25558);
  and AND_12231(g26394,g22530,g25560);
  and AND_12232(g26395,g22547,g25561);
  and AND_12233(g26397,g19475,g25563);
  and AND_12234(g26398,g24946,g10474);
  and AND_12235(g26399,g15572,g25566);
  and AND_12236(g26423,g19488,g24356);
  and AND_12237(g26484,g24946,g8841);
  and AND_12238(g26485,g24968,g10502);
  and AND_12239(g26486,g4423,g24358);
  and AND_12240(g26487,g15702,g24359);
  and AND_12241(g26511,g19265,g24364);
  and AND_12242(g26513,g19501,g24365);
  and AND_12243(g26514,g7400,g25564);
  and AND_12244(g26516,g24968,g8876);
  and AND_12245(g26517,g15708,g24367);
  and AND_12246(g26541,g319,g24375);
  and AND_12247(g26542,g13102,g24376);
  and AND_12248(g26543,g12910,g24377);
  and AND_12249(g26544,g7446,g24357);
  and AND_12250(g26547,g13283,g25027);
  and AND_12251(g26571,g10472,g24386);
  and AND_12252(g26572,g7443,g24439);
  and AND_12253(g26602,g7487,g24453);
  and AND_12254(g26604,g13248,g25051);
  and AND_12255(g26606,g1018,g24510);
  and AND_12256(g26610,g14198,g24405);
  and AND_12257(g26611,g24935,g20580);
  and AND_12258(g26612,g901,g24407);
  and AND_12259(g26613,g1361,g24518);
  and AND_12260(g26629,g14173,g24418);
  and AND_12261(g26630,g7592,g24419);
  and AND_12262(g26633,g24964,g20616);
  and AND_12263(g26635,g25321,g20617);
  and AND_12264(g26650,g10796,g24424);
  and AND_12265(g26651,g22707,g24425);
  and AND_12266(g26652,g10799,g24426);
  and AND_12267(g26670,g13385,g24428);
  and AND_12268(g26671,g316,g24429);
  and AND_12269(g26684,g25407,g20673);
  and AND_12270(g26689,g15754,g24431);
  and AND_12271(g26711,g25446,g20713);
  and AND_12272(g26712,g24508,g24463);
  and AND_12273(g26713,g25447,g20714);
  and AND_12274(g26719,g10709,g24438);
  and AND_12275(g26749,g24494,g23578);
  and AND_12276(g26750,g24514,g24474);
  and AND_12277(g26753,g16024,g24452);
  and AND_12278(g26778,g25501,g20923);
  and AND_12279(g26779,g24497,g23620);
  and AND_12280(g26780,g4098,g24437);
  and AND_12281(g26783,g25037,g21048);
  and AND_12282(g26799,g25247,g21068);
  and AND_12283(g26808,g25521,g21185);
  and AND_12284(g26815,g4108,g24528);
  and AND_12285(g26819,g106,g24490);
  and AND_12286(g26821,g24821,g13103);
  and AND_12287(g26822,g24841,g13116);
  and AND_12288(g26823,g24401,g13106);
  and AND_12289(g26826,g24907,g15747);
  and AND_12290(g26828,g24919,g15756);
  and AND_12291(g26829,g2844,g24505);
  and AND_12292(g26833,g2852,g24509);
  and AND_12293(g26838,g2860,g24515);
  and AND_12294(g26839,g2988,g24516);
  and AND_12295(g26842,g2894,g24522);
  and AND_12296(g26844,g25261,g21418);
  and AND_12297(g26845,g24391,g21426);
  and AND_12298(g26846,g37,g24524);
  and AND_12299(g26847,g2873,g24525);
  and AND_12300(g26848,g2950,g24526);
  and AND_12301(g26849,g2994,g24527);
  and AND_12302(g26852,g24975,g24958);
  and AND_12303(g26853,g94,g24533);
  and AND_12304(g26854,g2868,g24534);
  and AND_12305(g26855,g2960,g24535);
  and AND_12306(g26857,g25062,g25049);
  and AND_12307(g26858,g2970,g24540);
  and AND_12308(g26861,g25021,g25003);
  and AND_12309(g26863,g24974,g24957);
  and AND_12310(g26864,g2907,g24548);
  and AND_12311(g26871,g25038,g25020);
  and AND_12312(g26977,g23032,g26261,g26424,g25550);
  and AND_12313(g26994,g23032,g26226,g26424,g25557);
  and AND_12314(g27020,g4601,g25852);
  and AND_12315(g27025,g26334,g7917);
  and AND_12316(g27028,g26342,g1157);
  and AND_12317(g27029,g26327,g11031);
  and AND_12318(g27030,g26343,g7947);
  and AND_12319(g27032,g7704,g5180,g5188,g26200);
  and AND_12320(g27033,g25767,g19273);
  and AND_12321(g27034,g26328,g8609);
  and AND_12322(g27035,g26348,g1500);
  and AND_12323(g27036,g26329,g11038);
  and AND_12324(g27039,g7738,g5527,g5535,g26223);
  and AND_12325(g27040,g7812,g6565,g6573,g26226);
  and AND_12326(g27041,g8519,g26330);
  and AND_12327(g27042,g25774,g19343);
  and AND_12328(g27043,g26335,g8632);
  and AND_12329(g27044,g7766,g5873,g5881,g26241);
  and AND_12330(g27045,g10295,g3171,g3179,g26244);
  and AND_12331(g27050,g25789,g22338);
  and AND_12332(g27057,g7791,g6219,g6227,g26261);
  and AND_12333(g27058,g10323,g3522,g3530,g26264);
  and AND_12334(g27073,g7121,g3873,g3881,g26281);
  and AND_12335(g27083,g25819,g22456);
  and AND_12336(g27085,g25835,g22494);
  and AND_12337(g27086,g25836,g22495);
  and AND_12338(g27087,g13872,g26284);
  and AND_12339(g27090,g25997,g16423);
  and AND_12340(g27094,g25997,g16472);
  and AND_12341(g27095,g25997,g16473);
  and AND_12342(g27096,g26026,g16475);
  and AND_12343(g27097,g25867,g22526);
  and AND_12344(g27098,g25868,g22528);
  and AND_12345(g27099,g14094,g26352);
  and AND_12346(g27103,g25997,g16509);
  and AND_12347(g27104,g25997,g16510);
  and AND_12348(g27105,g26026,g16511);
  and AND_12349(g27106,g26026,g16512);
  and AND_12350(g27107,g26055,g16514);
  and AND_12351(g27113,g25997,g16522);
  and AND_12352(g27114,g25997,g16523);
  and AND_12353(g27115,g26026,g16526);
  and AND_12354(g27116,g26026,g16527);
  and AND_12355(g27117,g26055,g16528);
  and AND_12356(g27118,g26055,g16529);
  and AND_12357(g27119,g25877,g22542);
  and AND_12358(g27120,g25878,g22543);
  and AND_12359(g27121,g136,g26326);
  and AND_12360(g27127,g25997,g16582);
  and AND_12361(g27128,g25997,g16583);
  and AND_12362(g27129,g26026,g16584);
  and AND_12363(g27130,g26026,g16585);
  and AND_12364(g27131,g26055,g16588);
  and AND_12365(g27132,g26055,g16589);
  and AND_12366(g27134,g25997,g16602);
  and AND_12367(g27136,g26026,g16605);
  and AND_12368(g27137,g26026,g16606);
  and AND_12369(g27138,g26055,g16607);
  and AND_12370(g27139,g26055,g16608);
  and AND_12371(g27140,g25885,g22593);
  and AND_12372(g27145,g14121,g26382);
  and AND_12373(g27146,g26148,g8187,g1648);
  and AND_12374(g27148,g25997,g16622);
  and AND_12375(g27149,g25997,g16623);
  and AND_12376(g27151,g26026,g16626);
  and AND_12377(g27153,g26055,g16629);
  and AND_12378(g27154,g26055,g16630);
  and AND_12379(g27158,g26609,g16645);
  and AND_12380(g27160,g14163,g26340);
  and AND_12381(g27161,g26166,g8241,g1783);
  and AND_12382(g27162,g26171,g8259,g2208);
  and AND_12383(g27177,g25997,g16651);
  and AND_12384(g27178,g25997,g16652);
  and AND_12385(g27180,g26026,g16654);
  and AND_12386(g27181,g26026,g16655);
  and AND_12387(g27183,g26055,g16658);
  and AND_12388(g27184,g26628,g13756);
  and AND_12389(g27185,g26190,g8302,g1917);
  and AND_12390(g27186,g26195,g8316,g2342);
  and AND_12391(g27201,g25997,g16685);
  and AND_12392(g27202,g25997,g13876);
  and AND_12393(g27203,g26026,g16688);
  and AND_12394(g27204,g26026,g16689);
  and AND_12395(g27206,g26055,g16691);
  and AND_12396(g27207,g26055,g16692);
  and AND_12397(g27208,g9037,g26598);
  and AND_12398(g27209,g26213,g8365,g2051);
  and AND_12399(g27210,g26218,g8373,g2476);
  and AND_12400(g27211,g25997,g16716);
  and AND_12401(g27212,g25997,g16717);
  and AND_12402(g27213,g26026,g16721);
  and AND_12403(g27214,g26026,g13901);
  and AND_12404(g27215,g26055,g16724);
  and AND_12405(g27216,g26055,g16725);
  and AND_12406(g27217,g26236,g8418,g2610);
  and AND_12407(g27218,g25997,g16740);
  and AND_12408(g27219,g26026,g16742);
  and AND_12409(g27220,g26026,g16743);
  and AND_12410(g27221,g26055,g16747);
  and AND_12411(g27222,g26055,g13932);
  and AND_12412(g27227,g26026,g16771);
  and AND_12413(g27228,g26055,g16773);
  and AND_12414(g27229,g26055,g16774);
  and AND_12415(g27230,g25906,g19558);
  and AND_12416(g27234,g26055,g16814);
  and AND_12417(g27235,g25910,g19579);
  and AND_12418(g27246,g26690,g26673);
  and AND_12419(g27247,g2759,g26745);
  and AND_12420(g27249,g25929,g19678);
  and AND_12421(g27251,g26721,g26694);
  and AND_12422(g27252,g26733,g26703);
  and AND_12423(g27254,g25935,g19688);
  and AND_12424(g27255,g25936,g19689);
  and AND_12425(g27256,g25937,g19698);
  and AND_12426(g27259,g26755,g26725);
  and AND_12427(g27260,g26766,g26737);
  and AND_12428(g27262,g25997,g17092);
  and AND_12429(g27263,g25940,g19713);
  and AND_12430(g27264,g25941,g19714);
  and AND_12431(g27265,g26785,g26759);
  and AND_12432(g27266,g26789,g26770);
  and AND_12433(g27267,g26026,g17124);
  and AND_12434(g27268,g25942,g19733);
  and AND_12435(g27269,g25943,g19734);
  and AND_12436(g27270,g26805,g26793);
  and AND_12437(g27272,g26055,g17144);
  and AND_12438(g27275,g25945,g19745);
  and AND_12439(g27276,g9750,g26607);
  and AND_12440(g27277,g26359,g14191);
  and AND_12441(g27280,g9825,g26614);
  and AND_12442(g27281,g9830,g26615);
  and AND_12443(g27284,g9908,g26631);
  and AND_12444(g27285,g9912,g26632);
  and AND_12445(g27286,g6856,g26634);
  and AND_12446(g27287,g26545,g23011);
  and AND_12447(g27288,g26515,g23013);
  and AND_12448(g27291,g11969,g26653);
  and AND_12449(g27292,g1714,g26654);
  and AND_12450(g27293,g9972,g26655);
  and AND_12451(g27294,g9975,g26656);
  and AND_12452(g27298,g26573,g23026);
  and AND_12453(g27299,g26546,g23028);
  and AND_12454(g27300,g12370,g26672);
  and AND_12455(g27301,g11992,g26679);
  and AND_12456(g27302,g1848,g26680);
  and AND_12457(g27303,g11996,g26681);
  and AND_12458(g27304,g2273,g26682);
  and AND_12459(g27305,g10041,g26683);
  and AND_12460(g27309,g26603,g23057);
  and AND_12461(g27310,g26574,g23059);
  and AND_12462(g27311,g12431,g26693);
  and AND_12463(g27312,g12019,g26700);
  and AND_12464(g27313,g1982,g26701);
  and AND_12465(g27314,g12436,g26702);
  and AND_12466(g27315,g12022,g26709);
  and AND_12467(g27316,g2407,g26710);
  and AND_12468(g27323,g26268,g23086);
  and AND_12469(g27324,g10150,g26720);
  and AND_12470(g27325,g12478,g26724);
  and AND_12471(g27326,g12048,g26731);
  and AND_12472(g27327,g2116,g26732);
  and AND_12473(g27328,g12482,g26736);
  and AND_12474(g27329,g12052,g26743);
  and AND_12475(g27330,g2541,g26744);
  and AND_12476(g27331,g10177,g26754);
  and AND_12477(g27332,g12538,g26758);
  and AND_12478(g27333,g10180,g26765);
  and AND_12479(g27334,g12539,g26769);
  and AND_12480(g27335,g12087,g26776);
  and AND_12481(g27336,g2675,g26777);
  and AND_12482(g27339,g26400,g17308);
  and AND_12483(g27340,g10199,g26784);
  and AND_12484(g27341,g10203,g26788);
  and AND_12485(g27342,g12592,g26792);
  and AND_12486(g27346,g26400,g17389);
  and AND_12487(g27347,g26400,g17390);
  and AND_12488(g27348,g26488,g17392);
  and AND_12489(g27350,g10217,g26803);
  and AND_12490(g27351,g10218,g26804);
  and AND_12491(g27357,g26400,g17414);
  and AND_12492(g27358,g26400,g17415);
  and AND_12493(g27359,g26488,g17416);
  and AND_12494(g27360,g26488,g17417);
  and AND_12495(g27361,g26519,g17419);
  and AND_12496(g27362,g26080,g20036);
  and AND_12497(g27363,g10231,g26812);
  and AND_12498(g27369,g25894,g25324);
  and AND_12499(g27370,g26400,g17472);
  and AND_12500(g27371,g26400,g17473);
  and AND_12501(g27372,g26488,g17476);
  and AND_12502(g27373,g26488,g17477);
  and AND_12503(g27374,g26519,g17478);
  and AND_12504(g27375,g26519,g17479);
  and AND_12505(g27376,g26549,g17481);
  and AND_12506(g27378,g26089,g20052);
  and AND_12507(g27384,g26400,g17496);
  and AND_12508(g27385,g26400,g17497);
  and AND_12509(g27386,g26488,g17498);
  and AND_12510(g27387,g26488,g17499);
  and AND_12511(g27388,g26519,g17502);
  and AND_12512(g27389,g26519,g17503);
  and AND_12513(g27390,g26549,g17504);
  and AND_12514(g27391,g26549,g17505);
  and AND_12515(g27392,g26576,g17507);
  and AND_12516(g27393,g26099,g20066);
  and AND_12517(g27395,g8046,g26314,g9187,g9077);
  and AND_12518(g27404,g26400,g17518);
  and AND_12519(g27406,g26488,g17521);
  and AND_12520(g27407,g26488,g17522);
  and AND_12521(g27408,g26519,g17523);
  and AND_12522(g27409,g26519,g17524);
  and AND_12523(g27410,g26549,g17527);
  and AND_12524(g27411,g26549,g17528);
  and AND_12525(g27412,g26576,g17529);
  and AND_12526(g27413,g26576,g17530);
  and AND_12527(g27414,g255,g26827);
  and AND_12528(g27416,g8046,g26314,g9187,g504);
  and AND_12529(g27421,g8038,g26314,g9187,g9077);
  and AND_12530(g27427,g26400,g17575);
  and AND_12531(g27428,g26400,g17576);
  and AND_12532(g27430,g26488,g17579);
  and AND_12533(g27432,g26519,g17582);
  and AND_12534(g27433,g26519,g17583);
  and AND_12535(g27434,g26549,g17584);
  and AND_12536(g27435,g26549,g17585);
  and AND_12537(g27436,g26576,g17588);
  and AND_12538(g27437,g26576,g17589);
  and AND_12539(g27439,g232,g26831);
  and AND_12540(g27440,g8046,g26314,g518,g504);
  and AND_12541(g27445,g8038,g26314,g9187,g504);
  and AND_12542(g27451,g26400,g17599);
  and AND_12543(g27452,g26400,g17600);
  and AND_12544(g27454,g26488,g17602);
  and AND_12545(g27455,g26488,g17603);
  and AND_12546(g27457,g26519,g17606);
  and AND_12547(g27459,g26549,g17609);
  and AND_12548(g27460,g26549,g17610);
  and AND_12549(g27461,g26576,g17611);
  and AND_12550(g27462,g26576,g17612);
  and AND_12551(g27467,g269,g26832);
  and AND_12552(g27469,g8046,g26314,g518,g9077);
  and AND_12553(g27474,g8038,g26314,g518,g504);
  and AND_12554(g27480,g26400,g17638);
  and AND_12555(g27481,g26400,g14630);
  and AND_12556(g27482,g26488,g17641);
  and AND_12557(g27483,g26488,g17642);
  and AND_12558(g27485,g26519,g17644);
  and AND_12559(g27486,g26519,g17645);
  and AND_12560(g27488,g26549,g17648);
  and AND_12561(g27490,g26576,g17651);
  and AND_12562(g27491,g26576,g17652);
  and AND_12563(g27493,g246,g26837);
  and AND_12564(g27494,g8038,g26314,g518,g9077);
  and AND_12565(g27500,g26400,g17672);
  and AND_12566(g27501,g26400,g17673);
  and AND_12567(g27502,g26488,g17677);
  and AND_12568(g27503,g26488,g14668);
  and AND_12569(g27504,g26519,g17680);
  and AND_12570(g27505,g26519,g17681);
  and AND_12571(g27507,g26549,g17683);
  and AND_12572(g27508,g26549,g17684);
  and AND_12573(g27510,g26576,g17687);
  and AND_12574(g27517,g26400,g17707);
  and AND_12575(g27518,g26488,g17709);
  and AND_12576(g27519,g26488,g17710);
  and AND_12577(g27520,g26519,g17714);
  and AND_12578(g27521,g26519,g14700);
  and AND_12579(g27522,g26549,g17717);
  and AND_12580(g27523,g26549,g17718);
  and AND_12581(g27525,g26576,g17720);
  and AND_12582(g27526,g26576,g17721);
  and AND_12583(g27534,g26488,g17735);
  and AND_12584(g27535,g26519,g17737);
  and AND_12585(g27536,g26519,g17738);
  and AND_12586(g27537,g26549,g17742);
  and AND_12587(g27538,g26549,g14744);
  and AND_12588(g27539,g26576,g17745);
  and AND_12589(g27540,g26576,g17746);
  and AND_12590(g27541,g26278,g23334);
  and AND_12591(g27545,g26519,g17756);
  and AND_12592(g27546,g26549,g17758);
  and AND_12593(g27547,g26549,g17759);
  and AND_12594(g27548,g26576,g17763);
  and AND_12595(g27549,g26576,g14785);
  and AND_12596(g27553,g26293,g23353);
  and AND_12597(g27557,g26549,g17774);
  and AND_12598(g27558,g26576,g17776);
  and AND_12599(g27559,g26576,g17777);
  and AND_12600(g27560,g26299,g20191);
  and AND_12601(g27564,g26305,g23378);
  and AND_12602(g27568,g26576,g17791);
  and AND_12603(g27588,g26690,g26673);
  and AND_12604(g27594,g26721,g26694);
  and AND_12605(g27595,g26733,g26703);
  and AND_12606(g27598,g25899,g10475);
  and AND_12607(g27599,g26337,g20033);
  and AND_12608(g27600,g26755,g26725);
  and AND_12609(g27601,g26766,g26737);
  and AND_12610(g27602,g23032,g26244,g26424,g24966);
  and AND_12611(g27612,g25887,g8844);
  and AND_12612(g27614,g26785,g26759);
  and AND_12613(g27615,g26789,g26770);
  and AND_12614(g27616,g26349,g20449);
  and AND_12615(g27617,g23032,g26264,g26424,g24982);
  and AND_12616(g27627,g13266,g25790);
  and AND_12617(g27628,g26400,g18061);
  and AND_12618(g27633,g13076,g25766);
  and AND_12619(g27634,g26805,g26793);
  and AND_12620(g27635,g23032,g26281,g26424,g24996);
  and AND_12621(g27645,g26488,g15344);
  and AND_12622(g27646,g13094,g25773);
  and AND_12623(g27648,g25882,g8974);
  and AND_12624(g27649,g10820,g25820);
  and AND_12625(g27650,g26519,g15479);
  and AND_12626(g27651,g22448,g25781);
  and AND_12627(g27653,g26549,g15562);
  and AND_12628(g27658,g22491,g25786);
  and AND_12629(g27660,g24688,g26424,g22763);
  and AND_12630(g27661,g26576,g15568);
  and AND_12631(g27664,g1024,g25911);
  and AND_12632(g27665,g26872,g23519);
  and AND_12633(g27666,g26865,g23521);
  and AND_12634(g27667,g26361,g20601);
  and AND_12635(g27668,g1367,g25917);
  and AND_12636(g27669,g26840,g13278);
  and AND_12637(g27673,g25769,g23541);
  and AND_12638(g27674,g26873,g23543);
  and AND_12639(g27676,g26377,g20627);
  and AND_12640(g27677,g13021,g25888);
  and AND_12641(g27678,g947,g25830);
  and AND_12642(g27682,g25777,g23565);
  and AND_12643(g27683,g25770,g23567);
  and AND_12644(g27684,g26386,g20657);
  and AND_12645(g27685,g13032,g25895);
  and AND_12646(g27686,g1291,g25849);
  and AND_12647(g27690,g25784,g23607);
  and AND_12648(g27691,g25778,g23609);
  and AND_12649(g27692,g26392,g20697);
  and AND_12650(g27696,g25800,g23647);
  and AND_12651(g27697,g25785,g23649);
  and AND_12652(g27699,g26396,g20766);
  and AND_12653(g27700,g22342,g25182,g26424,g26148);
  and AND_12654(g27710,g26422,g20904);
  and AND_12655(g27711,g22369,g25193,g26424,g26166);
  and AND_12656(g27714,g22384,g25195,g26424,g26171);
  and AND_12657(g27723,g26512,g21049);
  and AND_12658(g27724,g22417,g25208,g26424,g26190);
  and AND_12659(g27727,g22432,g25211,g26424,g26195);
  and AND_12660(g27759,g22457,g25224,g26424,g26213);
  and AND_12661(g27762,g22472,g25226,g26424,g26218);
  and AND_12662(g27765,g4146,g25886);
  and AND_12663(g27817,g22498,g25245,g26424,g26236);
  and AND_12664(g27820,g7670,g25932);
  and AND_12665(g27821,g7680,g25892);
  and AND_12666(g27822,g4157,g25893);
  and AND_12667(g27932,g25944,g19369);
  and AND_12668(g27957,g25947,g15995);
  and AND_12669(g27958,g25950,g22449);
  and AND_12670(g27959,g25948,g19374);
  and AND_12671(g27962,g25954,g19597);
  and AND_12672(g27963,g25952,g16047);
  and AND_12673(g27964,g25956,g22492);
  and AND_12674(g27965,g25834,g13117);
  and AND_12675(g27968,g25958,g19614);
  and AND_12676(g27981,g26751,g23924);
  and AND_12677(g27988,g26781,g23941);
  and AND_12678(g27992,g26800,g23964);
  and AND_12679(g27995,g26809,g23985);
  and AND_12680(g27997,g26813,g23995);
  and AND_12681(g27999,g23032,g26200,g26424,g25529);
  and AND_12682(g28010,g23032,g26223,g26424,g25535);
  and AND_12683(g28020,g23032,g26241,g26424,g25542);
  and AND_12684(I26530,g26365,g24096,g24097,g24098);
  and AND_12685(I26531,g24099,g24100,g24101,g24102);
  and AND_12686(g28035,g24103,I26530,I26531);
  and AND_12687(g28107,g27970,g18874);
  and AND_12688(g28108,g7975,g27237);
  and AND_12689(g28110,g27974,g18886);
  and AND_12690(g28111,g27343,g22716);
  and AND_12691(g28112,g27352,g26162);
  and AND_12692(g28113,g8016,g27242);
  and AND_12693(g28114,g25869,g27051);
  and AND_12694(g28115,g27354,g22759);
  and AND_12695(g28116,g27366,g26183);
  and AND_12696(g28117,g8075,g27245);
  and AND_12697(g28124,g27368,g22842);
  and AND_12698(g28125,g27381,g26209);
  and AND_12699(g28130,g27353,g23063);
  and AND_12700(g28133,g27367,g23108);
  and AND_12701(g28136,g27382,g23135);
  and AND_12702(g28139,g27337,g26054);
  and AND_12703(g28141,g10831,g11797,g11261,g27163);
  and AND_12704(g28143,g27344,g26083);
  and AND_12705(g28144,g4608,g27020);
  and AND_12706(g28148,g27355,g26093);
  and AND_12707(g28150,g10862,g11834,g11283,g27187);
  and AND_12708(g28151,g8426,g27295);
  and AND_12709(g28152,g26297,g27279);
  and AND_12710(g28153,g26424,g22763,g27031);
  and AND_12711(g28154,g8492,g27306);
  and AND_12712(g28158,g26424,g22763,g27037);
  and AND_12713(g28159,g8553,g27317);
  and AND_12714(g28160,g26309,g27463);
  and AND_12715(g28164,g8651,g27528);
  and AND_12716(g28165,g27018,g22455);
  and AND_12717(g28171,g27016,g19385);
  and AND_12718(g28178,g27019,g19397);
  and AND_12719(g28182,g8770,g27349);
  and AND_12720(g28183,g27024,g19421);
  and AND_12721(g28185,g27026,g19435);
  and AND_12722(g28192,g8891,g27415);
  and AND_12723(g28193,g8851,g27629);
  and AND_12724(g28197,g27647,g11344);
  and AND_12725(g28198,g26649,g27492);
  and AND_12726(g28199,g27479,g16684);
  and AND_12727(g28200,g27652,g11383);
  and AND_12728(g28201,g27499,g16720);
  and AND_12729(g28202,g27659,g11413);
  and AND_12730(g28204,g26098,g27654);
  and AND_12731(g28205,g27516,g16746);
  and AND_12732(g28210,g9229,g27554);
  and AND_12733(g28213,g27720,g23380);
  and AND_12734(g28214,g27731,g26625);
  and AND_12735(g28215,g9264,g27565);
  and AND_12736(g28217,g27733,g23391);
  and AND_12737(g28218,g27768,g26645);
  and AND_12738(g28219,g9316,g27573);
  and AND_12739(g28223,g27338,g17194);
  and AND_12740(g28224,g27163,g22763,g27064);
  and AND_12741(g28225,g27770,g23400);
  and AND_12742(g28226,g27825,g26667);
  and AND_12743(g28227,g9397,g27583);
  and AND_12744(g28228,g27126,g19636);
  and AND_12745(g28229,g27345,g17213);
  and AND_12746(g28231,g27187,g22763,g27074);
  and AND_12747(g28232,g27732,g23586);
  and AND_12748(g28233,g27827,g23411);
  and AND_12749(g28234,g27877,g26686);
  and AND_12750(g28235,g9467,g27592);
  and AND_12751(g28236,g8515,g27971);
  and AND_12752(g28237,g9492,g27597);
  and AND_12753(g28238,g27133,g19658);
  and AND_12754(g28239,g27135,g19659);
  and AND_12755(g28240,g27356,g17239);
  and AND_12756(g28242,g27769,g23626);
  and AND_12757(g28243,g27879,g23423);
  and AND_12758(g28244,g27926,g26715);
  and AND_12759(g28245,g11367,g27975);
  and AND_12760(g28246,g8572,g27976);
  and AND_12761(g28247,g27147,g19675);
  and AND_12762(g28248,g27150,g19676);
  and AND_12763(g28249,g27152,g19677);
  and AND_12764(g28251,g27826,g23662);
  and AND_12765(g28252,g27159,g19682);
  and AND_12766(g28253,g23719,g27700);
  and AND_12767(g28254,g7268,g1668,g27395);
  and AND_12768(g28255,g8515,g27983);
  and AND_12769(g28256,g11398,g27984);
  and AND_12770(g28257,g27179,g19686);
  and AND_12771(g28258,g27182,g19687);
  and AND_12772(g28260,g27703,g26518);
  and AND_12773(g28261,g27878,g23695);
  and AND_12774(g28263,g23747,g27711);
  and AND_12775(g28264,g7315,g1802,g27416);
  and AND_12776(g28265,g11367,g27989);
  and AND_12777(g28266,g23748,g27714);
  and AND_12778(g28267,g7328,g2227,g27421);
  and AND_12779(g28268,g8572,g27990);
  and AND_12780(g28269,g27205,g19712);
  and AND_12781(g28272,g27721,g26548);
  and AND_12782(g28273,g27927,g23729);
  and AND_12783(g28280,g23761,g27724);
  and AND_12784(g28281,g7362,g1936,g27440);
  and AND_12785(g28282,g23762,g27727);
  and AND_12786(g28283,g7380,g2361,g27445);
  and AND_12787(g28284,g11398,g27994);
  and AND_12788(g28285,g9657,g27717);
  and AND_12789(g28289,g27734,g26575);
  and AND_12790(g28290,g23780,g27759);
  and AND_12791(g28291,g7411,g2070,g27469);
  and AND_12792(g28292,g23781,g27762);
  and AND_12793(g28293,g7424,g2495,g27474);
  and AND_12794(g28299,g9716,g27670);
  and AND_12795(g28300,g27771,g26605);
  and AND_12796(g28301,g27224,g19750);
  and AND_12797(g28302,g23809,g27817);
  and AND_12798(g28303,g7462,g2629,g27494);
  and AND_12799(g28304,g27226,g19753);
  and AND_12800(g28311,g9792,g27679);
  and AND_12801(g28312,g27828,g26608);
  and AND_12802(g28313,g27231,g19766);
  and AND_12803(g28314,g27552,g14205);
  and AND_12804(g28315,g27232,g19769);
  and AND_12805(g28318,g27233,g19770);
  and AND_12806(g28324,g9875,g27687);
  and AND_12807(g28327,g27365,g19785);
  and AND_12808(g28330,g27238,g19786);
  and AND_12809(g28333,g27239,g19787);
  and AND_12810(g28339,g9946,g27693);
  and AND_12811(g28341,g27240,g19790);
  and AND_12812(g28343,g27380,g19799);
  and AND_12813(g28346,g27243,g19800);
  and AND_12814(g28352,g10014,g27705);
  and AND_12815(g28360,g27401,g19861);
  and AND_12816(g28415,g27250,g19963);
  and AND_12817(g28426,g27257,g20006);
  and AND_12818(g28427,g27258,g20008);
  and AND_12819(g28439,g27273,g10233);
  and AND_12820(g28440,g27274,g20059);
  and AND_12821(g28442,g27278,g20072);
  and AND_12822(g28451,g27283,g20090);
  and AND_12823(g28453,g27582,g10233);
  and AND_12824(g28454,g26976,g12233);
  and AND_12825(g28455,g27289,g20103);
  and AND_12826(g28456,g27290,g20104);
  and AND_12827(I26948,g24981,g26424,g22698);
  and AND_12828(g28458,g27187,g12730,g20887,I26948);
  and AND_12829(g28466,g27960,g17637);
  and AND_12830(g28467,g26993,g12295);
  and AND_12831(I26960,g24995,g26424,g22698);
  and AND_12832(g28471,g27187,g12762,g21024,I26960);
  and AND_12833(g28477,g27966,g17676);
  and AND_12834(g28478,g27007,g12345);
  and AND_12835(I26972,g25011,g26424,g22698);
  and AND_12836(g28484,g27187,g10290,g21163,I26972);
  and AND_12837(g28488,g27969,g17713);
  and AND_12838(g28489,g27010,g12417);
  and AND_12839(g28494,g27973,g17741);
  and AND_12840(g28495,g27012,g12465);
  and AND_12841(g28499,g27982,g17762);
  and AND_12842(g28523,g27704,g15585);
  and AND_12843(g28524,g6821,g27084);
  and AND_12844(g28528,g27187,g12730);
  and AND_12845(g28530,g27383,g20240);
  and AND_12846(g28531,g27722,g15608);
  and AND_12847(g28532,g27394,g20265);
  and AND_12848(g28535,g11981,g27088);
  and AND_12849(g28537,g6832,g27089);
  and AND_12850(g28539,g27187,g12762);
  and AND_12851(g28541,g27403,g20274);
  and AND_12852(g28542,g27405,g20275);
  and AND_12853(g28543,g27735,g15628);
  and AND_12854(g28547,g6821,g27091);
  and AND_12855(g28550,g12009,g27092);
  and AND_12856(g28553,g27187,g10290);
  and AND_12857(g28554,g27426,g20372);
  and AND_12858(g28555,g27429,g20373);
  and AND_12859(g28556,g27431,g20374);
  and AND_12860(g28557,g27772,g15647);
  and AND_12861(g28558,g7301,g27046);
  and AND_12862(g28563,g11981,g27100);
  and AND_12863(g28567,g6832,g27101);
  and AND_12864(g28569,g27453,g20433);
  and AND_12865(g28570,g27456,g20434);
  and AND_12866(g28571,g27458,g20435);
  and AND_12867(g28572,g27829,g15669);
  and AND_12868(g28573,g7349,g27059);
  and AND_12869(g28583,g12009,g27112);
  and AND_12870(g28585,g27063,g10530);
  and AND_12871(g28586,g27484,g20497);
  and AND_12872(g28587,g27487,g20498);
  and AND_12873(g28588,g27489,g20499);
  and AND_12874(g28597,g27515,g20508);
  and AND_12875(g28599,g27027,g8922);
  and AND_12876(g28601,g27506,g20514);
  and AND_12877(g28602,g27509,g20515);
  and AND_12878(g28612,g27524,g20539);
  and AND_12879(g28616,g27532,g20551);
  and AND_12880(g28617,g27533,g20552);
  and AND_12881(g28624,g22357,g27009);
  and AND_12882(g28626,g27542,g20573);
  and AND_12883(g28627,g27543,g20574);
  and AND_12884(g28630,g27544,g20575);
  and AND_12885(g28637,g22399,g27011);
  and AND_12886(g28638,g27551,g20583);
  and AND_12887(g28639,g27767,g20597);
  and AND_12888(g28642,g27555,g20598);
  and AND_12889(g28645,g27556,g20599);
  and AND_12890(g28652,g27282,g10288);
  and AND_12891(g28653,g7544,g27014);
  and AND_12892(g28654,g1030,g27108);
  and AND_12893(g28655,g27561,g20603);
  and AND_12894(g28657,g27562,g20606);
  and AND_12895(g28658,g27563,g20611);
  and AND_12896(g28660,g27824,g20623);
  and AND_12897(g28663,g27566,g20624);
  and AND_12898(g28666,g27567,g20625);
  and AND_12899(g28672,g7577,g27017);
  and AND_12900(g28673,g1373,g27122);
  and AND_12901(g28674,g27569,g20629);
  and AND_12902(g28676,g27570,g20632);
  and AND_12903(g28677,g27571,g20635);
  and AND_12904(g28679,g27572,g20638);
  and AND_12905(g28683,g27876,g20649);
  and AND_12906(g28686,g27574,g20650);
  and AND_12907(g28689,g27575,g20651);
  and AND_12908(g28692,g27578,g20661);
  and AND_12909(g28694,g27579,g20664);
  and AND_12910(g28695,g27580,g20666);
  and AND_12911(g28697,g27581,g20669);
  and AND_12912(g28703,g27925,g20680);
  and AND_12913(g28706,g27584,g20681);
  and AND_12914(g28710,g27589,g20703);
  and AND_12915(g28712,g27590,g20708);
  and AND_12916(g28714,g27591,g20711);
  and AND_12917(g28722,g27955,g20738);
  and AND_12918(g28725,g27596,g20779);
  and AND_12919(g28739,g21434,g26424,g25274,g27395);
  and AND_12920(g28761,g21434,g26424,g25299,g27416);
  and AND_12921(g28768,g21434,g26424,g25308,g27421);
  and AND_12922(g28789,g21434,g26424,g25340,g27440);
  and AND_12923(g28799,g21434,g26424,g25348,g27445);
  and AND_12924(g28812,g26972,g13037);
  and AND_12925(g28813,g4104,g27038);
  and AND_12926(g28833,g21434,g26424,g25388,g27469);
  and AND_12927(g28846,g21434,g26424,g25399,g27474);
  and AND_12928(g28880,g21434,g26424,g25438,g27494);
  and AND_12929(g28889,g17292,g25169,g26424,g27395);
  and AND_12930(g28919,g27663,g21295);
  and AND_12931(g28924,g17317,g25183,g26424,g27416);
  and AND_12932(g28939,g17321,g25184,g26424,g27421);
  and AND_12933(g28959,g17401,g25194,g26424,g27440);
  and AND_12934(g28970,g17405,g25196,g26424,g27445);
  and AND_12935(I27349,g25534,g26424,g22698);
  and AND_12936(g28982,g27163,g12687,g20682,I27349);
  and AND_12937(g28991,g14438,g25209,g26424,g27469);
  and AND_12938(g28998,g17424,g25212,g26424,g27474);
  and AND_12939(I27364,g25541,g26424,g22698);
  and AND_12940(g29008,g27163,g12730,g20739,I27364);
  and AND_12941(g29029,g14506,g25227,g26424,g27494);
  and AND_12942(I27381,g25549,g26424,g22698);
  and AND_12943(g29036,g27163,g12762,g20875,I27381);
  and AND_12944(I27409,g25556,g26424,g22698);
  and AND_12945(g29073,g27163,g10290,g21012,I27409);
  and AND_12946(I27429,g25562,g26424,g22698);
  and AND_12947(g29110,g27187,g12687,g20751,I27429);
  and AND_12948(g29178,g27163,g12687);
  and AND_12949(g29182,g27163,g12730);
  and AND_12950(g29188,g27163,g12762);
  and AND_12951(g29192,g27163,g10290);
  and AND_12952(g29199,g27187,g12687);
  and AND_12953(I27503,g19890,g24075,g24076,g28032);
  and AND_12954(I27504,g24077,g24078,g24079,g24080);
  and AND_12955(g29201,g24081,I27503,I27504);
  and AND_12956(I27508,g19935,g24082,g24083,g28033);
  and AND_12957(I27509,g24084,g24085,g24086,g24087);
  and AND_12958(g29202,g24088,I27508,I27509);
  and AND_12959(I27513,g19984,g24089,g24090,g28034);
  and AND_12960(I27514,g24091,g24092,g24093,g24094);
  and AND_12961(g29203,g24095,I27513,I27514);
  and AND_12962(I27518,g20720,g24104,g24105,g24106);
  and AND_12963(I27519,g28036,g24107,g24108,g24109);
  and AND_12964(g29204,g24110,I27518,I27519);
  and AND_12965(I27523,g20857,g24111,g24112,g24113);
  and AND_12966(I27524,g28037,g24114,g24115,g24116);
  and AND_12967(g29205,g24117,I27523,I27524);
  and AND_12968(I27528,g20998,g24118,g24119,g24120);
  and AND_12969(I27529,g28038,g24121,g24122,g24123);
  and AND_12970(g29206,g24124,I27528,I27529);
  and AND_12971(I27533,g21143,g24125,g24126,g24127);
  and AND_12972(I27534,g28039,g24128,g24129,g24130);
  and AND_12973(g29207,g24131,I27533,I27534);
  and AND_12974(I27538,g21209,g24132,g24133,g24134);
  and AND_12975(I27539,g28040,g24135,g24136,g24137);
  and AND_12976(g29208,g24138,I27538,I27539);
  and AND_12977(g29314,g29005,g22144);
  and AND_12978(g29315,g29188,g7051,g5990);
  and AND_12979(g29316,g28528,g6875,g3288);
  and AND_12980(g29320,g29068,g22147);
  and AND_12981(g29321,g29033,g22148);
  and AND_12982(g29322,g29192,g7074,g6336);
  and AND_12983(g29323,g28539,g6905,g3639);
  and AND_12984(g29324,g29078,g18883);
  and AND_12985(g29326,g29105,g22155);
  and AND_12986(g29327,g29070,g22156);
  and AND_12987(g29328,g28553,g6928,g3990);
  and AND_12988(g29329,g7995,g28353);
  and AND_12989(g29330,g29114,g18894);
  and AND_12990(g29331,g29143,g22169);
  and AND_12991(g29332,g29107,g22170);
  and AND_12992(g29334,g29148,g18908);
  and AND_12993(g29336,g4704,g28363);
  and AND_12994(g29337,g29166,g22180);
  and AND_12995(g29338,g29145,g22181);
  and AND_12996(g29344,g29168,g18932);
  and AND_12997(g29345,g4749,g28376);
  and AND_12998(g29346,g4894,g28381);
  and AND_12999(g29347,g29176,g22201);
  and AND_13000(g29349,g4760,g28391);
  and AND_13001(g29350,g4939,g28395);
  and AND_13002(g29351,g4771,g28406);
  and AND_13003(g29352,g4950,g28410);
  and AND_13004(g29354,g4961,g28421);
  and AND_13005(g29360,g27364,g28294);
  and AND_13006(g29362,g27379,g28307);
  and AND_13007(g29363,g8458,g28444);
  and AND_13008(g29364,g27400,g28321);
  and AND_13009(g29367,g8575,g28325);
  and AND_13010(g29369,g28209,g22341);
  and AND_13011(g29375,g13946,g28370);
  and AND_13012(g29376,g14002,g28504);
  and AND_13013(g29377,g28132,g19387);
  and AND_13014(g29378,g28137,g22493);
  and AND_13015(g29380,g28134,g19396);
  and AND_13016(g29381,g28135,g19399);
  and AND_13017(g29382,g26424,g22763,g28172);
  and AND_13018(g29383,g28138,g19412);
  and AND_13019(g29384,g26424,g22763,g28179);
  and AND_13020(g29475,g14033,g28500);
  and AND_13021(g29477,g14090,g28441);
  and AND_13022(g29494,g9073,g28479);
  and AND_13023(g29509,g1600,g28755);
  and AND_13024(g29510,g28856,g22342);
  and AND_13025(g29511,g1736,g28783);
  and AND_13026(g29512,g2161,g28793);
  and AND_13027(g29513,g28448,g14095);
  and AND_13028(g29514,g1608,g28780);
  and AND_13029(g29515,g28888,g22342);
  and AND_13030(g29516,g28895,g22369);
  and AND_13031(g29517,g1870,g28827);
  and AND_13032(g29518,g28906,g22384);
  and AND_13033(g29519,g2295,g28840);
  and AND_13034(g29521,g1744,g28824);
  and AND_13035(g29522,g28923,g22369);
  and AND_13036(g29523,g28930,g22417);
  and AND_13037(g29524,g2004,g28864);
  and AND_13038(g29525,g2169,g28837);
  and AND_13039(g29526,g28938,g22384);
  and AND_13040(g29527,g28945,g22432);
  and AND_13041(g29528,g2429,g28874);
  and AND_13042(g29530,g1612,g28820);
  and AND_13043(g29531,g1664,g28559);
  and AND_13044(g29532,g1878,g28861);
  and AND_13045(g29533,g28958,g22417);
  and AND_13046(g29534,g28965,g22457);
  and AND_13047(g29535,g2303,g28871);
  and AND_13048(g29536,g28969,g22432);
  and AND_13049(g29537,g28976,g22472);
  and AND_13050(g29538,g2563,g28914);
  and AND_13051(g29547,g1748,g28857);
  and AND_13052(g29548,g1798,g28575);
  and AND_13053(g29549,g2012,g28900);
  and AND_13054(g29550,g28990,g22457);
  and AND_13055(g29551,g2173,g28867);
  and AND_13056(g29552,g2223,g28579);
  and AND_13057(g29553,g2437,g28911);
  and AND_13058(g29554,g28997,g22472);
  and AND_13059(g29555,g29004,g22498);
  and AND_13060(g29563,g1616,g28853);
  and AND_13061(g29564,g1882,g28896);
  and AND_13062(g29565,g1932,g28590);
  and AND_13063(g29566,g2307,g28907);
  and AND_13064(g29567,g2357,g28593);
  and AND_13065(g29568,g2571,g28950);
  and AND_13066(g29569,g29028,g22498);
  and AND_13067(g29570,g2763,g28598);
  and AND_13068(g29571,g28452,g11762);
  and AND_13069(g29572,g1620,g28885);
  and AND_13070(g29573,g1752,g28892);
  and AND_13071(g29574,g2016,g28931);
  and AND_13072(g29575,g2066,g28604);
  and AND_13073(g29576,g2177,g28903);
  and AND_13074(g29577,g2441,g28946);
  and AND_13075(g29578,g2491,g28606);
  and AND_13076(g29579,g28457,g7964);
  and AND_13077(g29580,g28519,g14186);
  and AND_13078(g29581,g28462,g11796);
  and AND_13079(g29582,g27766,g28608);
  and AND_13080(g29584,g1706,g29018);
  and AND_13081(g29585,g1756,g28920);
  and AND_13082(g29586,g1886,g28927);
  and AND_13083(g29587,g2181,g28935);
  and AND_13084(g29588,g2311,g28942);
  and AND_13085(g29589,g2575,g28977);
  and AND_13086(g29590,g2625,g28615);
  and AND_13087(g29591,g28552,g11346);
  and AND_13088(g29592,g28469,g11832);
  and AND_13089(g29593,g28470,g7985);
  and AND_13090(g29594,g28529,g14192);
  and AND_13091(g29595,g28475,g11833);
  and AND_13092(g29596,g27823,g28620);
  and AND_13093(g29598,g28823,g22342);
  and AND_13094(g29599,g1710,g29018);
  and AND_13095(g29600,g1840,g29049);
  and AND_13096(g29601,g1890,g28955);
  and AND_13097(g29602,g2020,g28962);
  and AND_13098(g29603,g2265,g29060);
  and AND_13099(g29604,g2315,g28966);
  and AND_13100(g29605,g2445,g28973);
  and AND_13101(g29606,g28480,g8011);
  and AND_13102(g29607,g28509,g14208);
  and AND_13103(g29608,g28568,g11385);
  and AND_13104(g29609,g28482,g11861);
  and AND_13105(g29610,g28483,g8026);
  and AND_13106(g29611,g28540,g14209);
  and AND_13107(g29612,g27875,g28633);
  and AND_13108(g29613,g28208,g19763);
  and AND_13109(g29614,g28860,g22369);
  and AND_13110(g29615,g1844,g29049);
  and AND_13111(g29616,g1974,g29085);
  and AND_13112(g29617,g2024,g28987);
  and AND_13113(g29618,g28870,g22384);
  and AND_13114(g29619,g2269,g29060);
  and AND_13115(g29620,g2399,g29097);
  and AND_13116(g29621,g2449,g28994);
  and AND_13117(g29622,g2579,g29001);
  and AND_13118(g29623,g28496,g11563);
  and AND_13119(g29624,g28491,g8070);
  and AND_13120(g29625,g28514,g14226);
  and AND_13121(g29626,g28584,g11415);
  and AND_13122(g29627,g28493,g11884);
  and AND_13123(g29628,g27924,g28648);
  and AND_13124(g29629,g28211,g19779);
  and AND_13125(g29630,g28212,g19781);
  and AND_13126(g29631,g1682,g28656);
  and AND_13127(g29632,g28899,g22417);
  and AND_13128(g29633,g1978,g29085);
  and AND_13129(g29634,g2108,g29121);
  and AND_13130(g29635,g28910,g22432);
  and AND_13131(g29636,g2403,g29097);
  and AND_13132(g29637,g2533,g29134);
  and AND_13133(g29638,g2583,g29025);
  and AND_13134(g29639,g28510,g11618);
  and AND_13135(g29640,g28498,g8125);
  and AND_13136(g29641,g28520,g14237);
  and AND_13137(g29642,g27954,g28669);
  and AND_13138(g29644,g28216,g19794);
  and AND_13139(g29645,g1714,g29018);
  and AND_13140(g29646,g1816,g28675);
  and AND_13141(g29647,g28934,g22457);
  and AND_13142(g29648,g2112,g29121);
  and AND_13143(g29649,g2241,g28678);
  and AND_13144(g29650,g28949,g22472);
  and AND_13145(g29651,g2537,g29134);
  and AND_13146(g29652,g2667,g29157);
  and AND_13147(g29656,g28515,g11666);
  and AND_13148(g29661,g1687,g29015);
  and AND_13149(g29662,g1848,g29049);
  and AND_13150(g29663,g1950,g28693);
  and AND_13151(g29664,g2273,g29060);
  and AND_13152(g29665,g2375,g28696);
  and AND_13153(g29666,g28980,g22498);
  and AND_13154(g29667,g2671,g29157);
  and AND_13155(g29668,g28527,g14255);
  and AND_13156(g29683,g1821,g29046);
  and AND_13157(g29684,g1982,g29085);
  and AND_13158(g29685,g2084,g28711);
  and AND_13159(g29686,g2246,g29057);
  and AND_13160(g29687,g2407,g29097);
  and AND_13161(g29688,g2509,g28713);
  and AND_13162(g29693,g28207,g10233);
  and AND_13163(g29708,g1955,g29082);
  and AND_13164(g29709,g2116,g29121);
  and AND_13165(g29710,g2380,g29094);
  and AND_13166(g29711,g2541,g29134);
  and AND_13167(g29712,g2643,g28726);
  and AND_13168(g29718,g28512,g11136);
  and AND_13169(g29731,g2089,g29118);
  and AND_13170(g29732,g2514,g29131);
  and AND_13171(g29733,g2675,g29157);
  and AND_13172(g29736,g28522,g10233);
  and AND_13173(g29740,g2648,g29154);
  and AND_13174(g29742,g28288,g10233);
  and AND_13175(g29743,g28206,g10233);
  and AND_13176(g29746,g28279,g20037);
  and AND_13177(g29747,g28286,g23196);
  and AND_13178(g29749,g28295,g23214);
  and AND_13179(g29750,g28296,g23215);
  and AND_13180(g29751,g28297,g23216);
  and AND_13181(g29752,g28516,g10233);
  and AND_13182(g29757,g28305,g23221);
  and AND_13183(g29758,g28306,g23222);
  and AND_13184(g29759,g28308,g23226);
  and AND_13185(g29760,g28309,g23227);
  and AND_13186(g29761,g28310,g23228);
  and AND_13187(g29762,g28298,g10233);
  and AND_13188(g29766,g28316,g23235);
  and AND_13189(g29767,g28317,g23236);
  and AND_13190(g29769,g28319,g23237);
  and AND_13191(g29770,g28320,g23238);
  and AND_13192(g29771,g28322,g23242);
  and AND_13193(g29772,g28323,g23243);
  and AND_13194(g29773,g28203,g10233);
  and AND_13195(g29774,g28287,g10233);
  and AND_13196(g29782,g28328,g23245);
  and AND_13197(g29783,g28329,g23246);
  and AND_13198(g29784,g28331,g23247);
  and AND_13199(g29785,g28332,g23248);
  and AND_13200(g29787,g28334,g23249);
  and AND_13201(g29788,g28335,g23250);
  and AND_13202(g29789,g28270,g10233);
  and AND_13203(g29794,g28342,g23256);
  and AND_13204(g29795,g28344,g23257);
  and AND_13205(g29796,g28345,g23258);
  and AND_13206(g29797,g28347,g23259);
  and AND_13207(g29798,g28348,g23260);
  and AND_13208(g29799,g28271,g10233);
  and AND_13209(g29803,g28414,g26836);
  and AND_13210(g29804,g1592,g29014);
  and AND_13211(g29805,g28357,g23270);
  and AND_13212(g29806,g28358,g23271);
  and AND_13213(g29807,g28359,g23272);
  and AND_13214(g29808,g28361,g23273);
  and AND_13215(g29809,g28362,g23274);
  and AND_13216(g29810,g28259,g11317);
  and AND_13217(g29834,g28368,g23278);
  and AND_13218(g29835,g28326,g24866);
  and AND_13219(g29836,g28425,g26841);
  and AND_13220(g29837,g28369,g20144);
  and AND_13221(g29838,g1636,g29044);
  and AND_13222(g29839,g1728,g29045);
  and AND_13223(g29840,g2153,g29056);
  and AND_13224(g29841,g28371,g23283);
  and AND_13225(g29842,g28372,g23284);
  and AND_13226(g29843,g28373,g23289);
  and AND_13227(g29844,g28374,g23290);
  and AND_13228(g29845,g28375,g23291);
  and AND_13229(g29850,g28340,g24893);
  and AND_13230(g29851,g1668,g29079);
  and AND_13231(g29852,g1772,g29080);
  and AND_13232(g29853,g1862,g29081);
  and AND_13233(g29854,g2197,g29092);
  and AND_13234(g29855,g2287,g29093);
  and AND_13235(g29856,g28385,g23303);
  and AND_13236(g29857,g28386,g23304);
  and AND_13237(g29858,g28387,g23306);
  and AND_13238(g29859,g28388,g23307);
  and AND_13239(g29860,g28389,g23312);
  and AND_13240(g29861,g28390,g23313);
  and AND_13241(g29865,g1802,g29115);
  and AND_13242(g29866,g1906,g29116);
  and AND_13243(g29867,g1996,g29117);
  and AND_13244(g29868,g2227,g29128);
  and AND_13245(g29869,g2331,g29129);
  and AND_13246(g29870,g2421,g29130);
  and AND_13247(g29871,g28400,g23332);
  and AND_13248(g29872,g28401,g23333);
  and AND_13249(g29874,g28402,g23336);
  and AND_13250(g29875,g28403,g23337);
  and AND_13251(g29876,g28404,g23339);
  and AND_13252(g29877,g28405,g23340);
  and AND_13253(g29880,g1936,g29149);
  and AND_13254(g29881,g2040,g29150);
  and AND_13255(g29882,g2361,g29151);
  and AND_13256(g29883,g2465,g29152);
  and AND_13257(g29884,g2555,g29153);
  and AND_13258(g29885,g28416,g23350);
  and AND_13259(g29887,g28417,g23351);
  and AND_13260(g29888,g28418,g23352);
  and AND_13261(g29890,g28419,g23355);
  and AND_13262(g29891,g28420,g23356);
  and AND_13263(g29894,g2070,g29169);
  and AND_13264(g29895,g2495,g29170);
  and AND_13265(g29896,g2599,g29171);
  and AND_13266(g29899,g28428,g23375);
  and AND_13267(g29901,g28429,g23376);
  and AND_13268(g29902,g28430,g23377);
  and AND_13269(g29907,g2629,g29177);
  and AND_13270(g29909,g28435,g23388);
  and AND_13271(g29924,g13031,g29190);
  and AND_13272(g29926,g1604,g28736);
  and AND_13273(g29937,g13044,g29196);
  and AND_13274(g29938,g23552,g28889);
  and AND_13275(g29940,g1740,g28758);
  and AND_13276(g29943,g2165,g28765);
  and AND_13277(g29949,g23575,g28924);
  and AND_13278(g29951,g1874,g28786);
  and AND_13279(g29952,g23576,g28939);
  and AND_13280(g29954,g2299,g28796);
  and AND_13281(g29959,g28953,g12823);
  and AND_13282(g29962,g23616,g28959);
  and AND_13283(g29964,g2008,g28830);
  and AND_13284(g29966,g23617,g28970);
  and AND_13285(g29968,g2433,g28843);
  and AND_13286(g29969,g28121,g20509);
  and AND_13287(g29973,g28981,g9206);
  and AND_13288(g29974,g29173,g12914);
  and AND_13289(g29975,g28986,g10420);
  and AND_13290(g29979,g23655,g28991);
  and AND_13291(g29982,g23656,g28998);
  and AND_13292(g29984,g2567,g28877);
  and AND_13293(g29985,g28127,g20532);
  and AND_13294(g29986,g28468,g23473);
  and AND_13295(g29987,g29197,g26424,g22763);
  and AND_13296(g29988,g29187,g12235);
  and AND_13297(g29989,g29006,g10489);
  and AND_13298(g29990,g29007,g9239);
  and AND_13299(g29991,g29179,g12922);
  and AND_13300(g29992,g29012,g10490);
  and AND_13301(g30000,g23685,g29029);
  and AND_13302(g30001,g28490,g23486);
  and AND_13303(g30002,g28481,g23487);
  and AND_13304(g30003,g28149,g9021);
  and AND_13305(g30004,g28521,g25837);
  and AND_13306(g30005,g28230,g24394);
  and AND_13307(g30006,g29032,g9259);
  and AND_13308(g30007,g29141,g12929);
  and AND_13309(g30008,g29191,g12297);
  and AND_13310(g30009,g29034,g10518);
  and AND_13311(g30010,g29035,g9274);
  and AND_13312(g30011,g29183,g12930);
  and AND_13313(g30015,g29040,g10519);
  and AND_13314(g30023,g28508,g20570);
  and AND_13315(g30024,g28497,g23501);
  and AND_13316(g30025,g28492,g23502);
  and AND_13317(g30026,g28476,g25064);
  and AND_13318(g30027,g29104,g12550);
  and AND_13319(g30028,g29069,g9311);
  and AND_13320(g30029,g29164,g12936);
  and AND_13321(g30030,g29198,g12347);
  and AND_13322(g30031,g29071,g10540);
  and AND_13323(g30032,g29072,g9326);
  and AND_13324(g30033,g29189,g12937);
  and AND_13325(g30034,g29077,g10541);
  and AND_13326(g30035,g22539,g28120);
  and AND_13327(g30041,g28511,g23518);
  and AND_13328(g30042,g29142,g12601);
  and AND_13329(g30043,g29106,g9392);
  and AND_13330(g30044,g29174,g12944);
  and AND_13331(g30045,g29200,g12419);
  and AND_13332(g30046,g29108,g10564);
  and AND_13333(g30047,g29109,g9407);
  and AND_13334(g30048,g29193,g12945);
  and AND_13335(g30049,g13114,g28167);
  and AND_13336(g30050,g22545,g28126);
  and AND_13337(g30051,g28513,g20604);
  and AND_13338(g30056,g29165,g12659);
  and AND_13339(g30057,g29144,g9462);
  and AND_13340(g30058,g29180,g12950);
  and AND_13341(g30059,g28106,g12467);
  and AND_13342(g30060,g29146,g10581);
  and AND_13343(g30061,g1036,g28188);
  and AND_13344(g30062,g13129,g28174);
  and AND_13345(g30064,g28517,g20630);
  and AND_13346(g30066,g28518,g20636);
  and AND_13347(g30069,g29175,g12708);
  and AND_13348(g30070,g29167,g9529);
  and AND_13349(g30071,g29184,g12975);
  and AND_13350(g30073,g1379,g28194);
  and AND_13351(g30075,g28525,g20662);
  and AND_13352(g30078,g28526,g20667);
  and AND_13353(g30080,g28121,g20674);
  and AND_13354(g30082,g29181,g12752);
  and AND_13355(g30083,g28533,g20698);
  and AND_13356(g30084,g28534,g20700);
  and AND_13357(g30086,g28536,g20704);
  and AND_13358(g30089,g28538,g20709);
  and AND_13359(g30091,g28127,g20716);
  and AND_13360(g30094,g28544,g20767);
  and AND_13361(g30095,g28545,g20768);
  and AND_13362(g30096,g28546,g20770);
  and AND_13363(g30098,g28548,g20774);
  and AND_13364(g30099,g28549,g20776);
  and AND_13365(g30101,g28551,g20780);
  and AND_13366(g30107,g28560,g20909);
  and AND_13367(g30108,g28561,g20910);
  and AND_13368(g30109,g28562,g20912);
  and AND_13369(g30110,g28564,g20916);
  and AND_13370(g30111,g28565,g20917);
  and AND_13371(g30112,g28566,g20919);
  and AND_13372(g30118,g28574,g21050);
  and AND_13373(g30120,g28576,g21051);
  and AND_13374(g30121,g28577,g21052);
  and AND_13375(g30122,g28578,g21054);
  and AND_13376(g30124,g28580,g21055);
  and AND_13377(g30125,g28581,g21056);
  and AND_13378(g30126,g28582,g21058);
  and AND_13379(g30131,g28589,g21178);
  and AND_13380(g30133,g28591,g21179);
  and AND_13381(g30135,g28592,g21180);
  and AND_13382(g30137,g28594,g21181);
  and AND_13383(g30138,g28595,g21182);
  and AND_13384(g30139,g28596,g21184);
  and AND_13385(g30140,g28600,g23749);
  and AND_13386(g30145,g28603,g21247);
  and AND_13387(g30149,g28605,g21248);
  and AND_13388(g30151,g28607,g21249);
  and AND_13389(g30152,g28609,g23767);
  and AND_13390(g30153,g28610,g23768);
  and AND_13391(g30154,g28611,g23769);
  and AND_13392(g30158,g28613,g21274);
  and AND_13393(g30161,g28614,g21275);
  and AND_13394(g30164,g28618,g23787);
  and AND_13395(g30165,g28619,g23788);
  and AND_13396(g30166,g28621,g23792);
  and AND_13397(g30167,g28622,g23793);
  and AND_13398(g30168,g28623,g23794);
  and AND_13399(g30172,g28625,g21286);
  and AND_13400(g30173,g28118,g13082);
  and AND_13401(g30174,g28628,g23812);
  and AND_13402(g30175,g28629,g23813);
  and AND_13403(g30177,g28631,g23814);
  and AND_13404(g30178,g28632,g23815);
  and AND_13405(g30179,g28634,g23819);
  and AND_13406(g30180,g28635,g23820);
  and AND_13407(g30181,g28636,g23821);
  and AND_13408(g30185,g28640,g23838);
  and AND_13409(g30186,g28641,g23839);
  and AND_13410(g30187,g28643,g23840);
  and AND_13411(g30188,g28644,g23841);
  and AND_13412(g30190,g28646,g23842);
  and AND_13413(g30191,g28647,g23843);
  and AND_13414(g30192,g28649,g23847);
  and AND_13415(g30193,g28650,g23848);
  and AND_13416(g30194,g28651,g23849);
  and AND_13417(g30196,g28659,g23858);
  and AND_13418(g30197,g28661,g23859);
  and AND_13419(g30198,g28662,g23860);
  and AND_13420(g30199,g28664,g23861);
  and AND_13421(g30200,g28665,g23862);
  and AND_13422(g30202,g28667,g23863);
  and AND_13423(g30203,g28668,g23864);
  and AND_13424(g30204,g28670,g23868);
  and AND_13425(g30205,g28671,g23869);
  and AND_13426(g30207,g28680,g23874);
  and AND_13427(g30208,g28681,g23875);
  and AND_13428(g30209,g28682,g23876);
  and AND_13429(g30210,g28684,g23877);
  and AND_13430(g30211,g28685,g23878);
  and AND_13431(g30212,g28687,g23879);
  and AND_13432(g30213,g28688,g23880);
  and AND_13433(g30215,g28690,g23881);
  and AND_13434(g30216,g28691,g23882);
  and AND_13435(g30219,g28698,g23887);
  and AND_13436(g30220,g28699,g23888);
  and AND_13437(g30221,g28700,g23893);
  and AND_13438(g30222,g28701,g23894);
  and AND_13439(g30223,g28702,g23895);
  and AND_13440(g30224,g28704,g23896);
  and AND_13441(g30225,g28705,g23897);
  and AND_13442(g30226,g28707,g23898);
  and AND_13443(g30227,g28708,g23899);
  and AND_13444(g30228,g28715,g23903);
  and AND_13445(g30229,g28716,g23904);
  and AND_13446(g30230,g28717,g23906);
  and AND_13447(g30231,g28718,g23907);
  and AND_13448(g30232,g28719,g23912);
  and AND_13449(g30233,g28720,g23913);
  and AND_13450(g30234,g28721,g23914);
  and AND_13451(g30235,g28723,g23915);
  and AND_13452(g30236,g28724,g23916);
  and AND_13453(g30238,g28727,g23922);
  and AND_13454(g30239,g28728,g23923);
  and AND_13455(g30241,g28729,g23926);
  and AND_13456(g30242,g28730,g23927);
  and AND_13457(g30243,g28731,g23929);
  and AND_13458(g30244,g28732,g23930);
  and AND_13459(g30245,g28733,g23935);
  and AND_13460(g30246,g28734,g23936);
  and AND_13461(g30247,g28735,g23937);
  and AND_13462(g30248,g28743,g23938);
  and AND_13463(g30250,g28744,g23939);
  and AND_13464(g30251,g28745,g23940);
  and AND_13465(g30253,g28746,g23943);
  and AND_13466(g30254,g28747,g23944);
  and AND_13467(g30255,g28748,g23946);
  and AND_13468(g30256,g28749,g23947);
  and AND_13469(g30257,g28750,g23952);
  and AND_13470(g30258,g28751,g23953);
  and AND_13471(g30261,g28772,g23961);
  and AND_13472(g30263,g28773,g23962);
  and AND_13473(g30264,g28774,g23963);
  and AND_13474(g30266,g28775,g23966);
  and AND_13475(g30267,g28776,g23967);
  and AND_13476(g30268,g28777,g23969);
  and AND_13477(g30269,g28778,g23970);
  and AND_13478(g30272,g28814,g23982);
  and AND_13479(g30274,g28815,g23983);
  and AND_13480(g30275,g28816,g23984);
  and AND_13481(g30277,g28817,g23987);
  and AND_13482(g30278,g28818,g23988);
  and AND_13483(g30281,g28850,g23992);
  and AND_13484(g30283,g28851,g23993);
  and AND_13485(g30284,g28852,g23994);
  and AND_13486(g30289,g28884,g24000);
  and AND_13487(g30308,g29178,g7004,g5297);
  and AND_13488(g30315,g29182,g7028,g5644);
  and AND_13489(g30316,g29199,g7097,g6682);
  and AND_13490(g30564,g21358,g29385);
  and AND_13491(g30566,g26247,g29507);
  and AND_13492(g30576,g18898,g29800);
  and AND_13493(g30577,g26267,g29679);
  and AND_13494(g30583,g19666,g29355);
  and AND_13495(g30589,g18898,g29811);
  and AND_13496(g30590,g18911,g29812);
  and AND_13497(g30592,g30270,g18929);
  and AND_13498(g30594,g18898,g29846);
  and AND_13499(g30595,g18911,g29847);
  and AND_13500(g30596,g30279,g18947);
  and AND_13501(g30598,g18898,g29862);
  and AND_13502(g30599,g18911,g29863);
  and AND_13503(g30600,g30287,g18975);
  and AND_13504(g30604,g18911,g29878);
  and AND_13505(g30607,g30291,g18989);
  and AND_13506(g30612,g26338,g29597);
  and AND_13507(g30614,g20154,g29814);
  and AND_13508(g30670,g11330,g29359);
  and AND_13509(g30671,g29319,g22317);
  and AND_13510(g30673,g20175,g29814);
  and AND_13511(g30730,g26346,g29778);
  and AND_13512(g30731,g11374,g29361);
  and AND_13513(g30735,g29814,g22319);
  and AND_13514(g30825,g29814,g22332);
  and AND_13515(g30914,g29873,g20887);
  and AND_13516(g30915,g29886,g24778);
  and AND_13517(g30918,g8681,g29707);
  and AND_13518(g30919,g29898,g23286);
  and AND_13519(g30920,g29889,g21024);
  and AND_13520(g30921,g29900,g24789);
  and AND_13521(g30925,g29908,g23309);
  and AND_13522(g30926,g29903,g21163);
  and AND_13523(g30927,g29910,g24795);
  and AND_13524(g30930,g29915,g23342);
  and AND_13525(g30935,g8808,g29745);
  and AND_13526(g30936,g8830,g29916);
  and AND_13527(g30937,g22626,g29814);
  and AND_13528(g30982,g8895,g29933);
  and AND_13529(g31015,g29476,g22758);
  and AND_13530(g31016,g29478,g22840);
  and AND_13531(g31017,g29479,g22841);
  and AND_13532(g31018,g29480,g22855);
  and AND_13533(g31019,g29481,g22856);
  and AND_13534(g31021,g26025,g29814);
  and AND_13535(g31066,g29483,g22865);
  and AND_13536(g31067,g29484,g22868);
  and AND_13537(g31069,g29793,g14150);
  and AND_13538(g31070,g29814,g25985);
  and AND_13539(g31115,g29487,g22882);
  and AND_13540(g31118,g29490,g22906);
  and AND_13541(g31120,g1700,g29976);
  and AND_13542(g31122,g12144,g29993);
  and AND_13543(g31123,g1834,g29994);
  and AND_13544(g31124,g2259,g29997);
  and AND_13545(g31125,g29502,g22973);
  and AND_13546(g31128,g12187,g30016);
  and AND_13547(g31129,g1968,g30017);
  and AND_13548(g31130,g12191,g30019);
  and AND_13549(g31131,g2393,g30020);
  and AND_13550(g31132,g29504,g22987);
  and AND_13551(g31139,g12221,g30036);
  and AND_13552(g31140,g2102,g30037);
  and AND_13553(g31141,g12224,g30038);
  and AND_13554(g31142,g2527,g30039);
  and AND_13555(g31143,g29506,g22999);
  and AND_13556(g31145,g9970,g30052);
  and AND_13557(g31146,g12285,g30053);
  and AND_13558(g31147,g12286,g30054);
  and AND_13559(g31148,g2661,g30055);
  and AND_13560(g31149,g29508,g23021);
  and AND_13561(g31150,g1682,g30063);
  and AND_13562(g31151,g10037,g30065);
  and AND_13563(g31152,g10039,g30067);
  and AND_13564(g31153,g12336,g30068);
  and AND_13565(g31154,g19128,g29814);
  and AND_13566(g31166,g1816,g30074);
  and AND_13567(g31167,g10080,g30076);
  and AND_13568(g31168,g2241,g30077);
  and AND_13569(g31169,g10083,g30079);
  and AND_13570(g31170,g19128,g29814);
  and AND_13571(g31182,g30240,g20682);
  and AND_13572(g31183,g30249,g25174);
  and AND_13573(g31184,g1950,g30085);
  and AND_13574(g31185,g10114,g30087);
  and AND_13575(g31186,g2375,g30088);
  and AND_13576(g31187,g10118,g30090);
  and AND_13577(g31188,g20028,g29653);
  and AND_13578(g31194,g19128,g29814);
  and AND_13579(g31206,g30260,g23890);
  and AND_13580(g31207,g30252,g20739);
  and AND_13581(g31208,g30262,g25188);
  and AND_13582(g31209,g2084,g30097);
  and AND_13583(g31210,g2509,g30100);
  and AND_13584(g31211,g10156,g30102);
  and AND_13585(g31212,g20028,g29669);
  and AND_13586(g31218,g30271,g23909);
  and AND_13587(g31219,g30265,g20875);
  and AND_13588(g31220,g30273,g25202);
  and AND_13589(g31222,g2643,g30113);
  and AND_13590(g31223,g20028,g29689);
  and AND_13591(g31224,g30280,g23932);
  and AND_13592(g31225,g30276,g21012);
  and AND_13593(g31226,g30282,g25218);
  and AND_13594(g31228,g20028,g29713);
  and AND_13595(g31229,g30288,g23949);
  and AND_13596(g31230,g30285,g20751);
  and AND_13597(g31231,g30290,g25239);
  and AND_13598(g31232,g30294,g23972);
  and AND_13599(g31237,g29366,g25325);
  and AND_13600(g31238,g29583,g20053);
  and AND_13601(g31240,g14793,g30206);
  and AND_13602(g31242,g29373,g25409);
  and AND_13603(g31252,g29643,g20101);
  and AND_13604(g31261,g14754,g30259);
  and AND_13605(g31266,g30129,g27742);
  and AND_13606(g31270,g29692,g23282);
  and AND_13607(g31271,g29706,g23300);
  and AND_13608(g31272,g30117,g27742);
  and AND_13609(g31273,g30143,g27779);
  and AND_13610(g31275,g30147,g27800);
  and AND_13611(g31278,g29716,g23302);
  and AND_13612(g31280,g29717,g23305);
  and AND_13613(g31281,g30106,g27742);
  and AND_13614(g31282,g30130,g27779);
  and AND_13615(g31283,g30156,g27837);
  and AND_13616(g31285,g30134,g27800);
  and AND_13617(g31286,g30159,g27858);
  and AND_13618(g31290,g29734,g23335);
  and AND_13619(g31292,g29735,g23338);
  and AND_13620(g31296,g30119,g27779);
  and AND_13621(g31297,g30144,g27837);
  and AND_13622(g31298,g30169,g27886);
  and AND_13623(g31299,g30123,g27800);
  and AND_13624(g31300,g30148,g27858);
  and AND_13625(g31301,g30170,g27907);
  and AND_13626(g31305,g29741,g23354);
  and AND_13627(g31309,g30132,g27837);
  and AND_13628(g31310,g30157,g27886);
  and AND_13629(g31312,g30136,g27858);
  and AND_13630(g31313,g30160,g27907);
  and AND_13631(g31314,g30183,g27937);
  and AND_13632(g31321,g30146,g27886);
  and AND_13633(g31323,g30150,g27907);
  and AND_13634(g31324,g30171,g27937);
  and AND_13635(g31327,g19200,g29814);
  and AND_13636(g31374,g29748,g23390);
  and AND_13637(g31376,g24952,g29814);
  and AND_13638(g31467,g30162,g27937);
  and AND_13639(g31470,g29753,g23398);
  and AND_13640(g31471,g29754,g23399);
  and AND_13641(g31475,g29756,g23406);
  and AND_13642(g31477,g29763,g23409);
  and AND_13643(g31478,g29764,g23410);
  and AND_13644(g31480,g1644,g30296);
  and AND_13645(g31481,g29768,g23417);
  and AND_13646(g31484,g29775,g23418);
  and AND_13647(g31485,g29776,g23421);
  and AND_13648(g31486,g29777,g23422);
  and AND_13649(g31488,g1779,g30302);
  and AND_13650(g31489,g2204,g30305);
  and AND_13651(g31490,g29786,g23429);
  and AND_13652(g31492,g29790,g23431);
  and AND_13653(g31493,g29791,g23434);
  and AND_13654(g31494,g29792,g23435);
  and AND_13655(g31495,g1913,g30309);
  and AND_13656(g31496,g2338,g30312);
  and AND_13657(g31497,g20041,g29930);
  and AND_13658(g31499,g29801,g23446);
  and AND_13659(g31500,g29802,g23449);
  and AND_13660(g31501,g2047,g29310);
  and AND_13661(g31502,g2472,g29311);
  and AND_13662(g31503,g20041,g29945);
  and AND_13663(g31504,g29370,g10553);
  and AND_13664(g31505,g30195,g24379);
  and AND_13665(g31508,g29813,g23459);
  and AND_13666(g31513,g2606,g29318);
  and AND_13667(g31514,g20041,g29956);
  and AND_13668(g31516,g29848,g23476);
  and AND_13669(g31517,g29849,g23482);
  and AND_13670(g31518,g20041,g29970);
  and AND_13671(g31519,g29864,g23490);
  and AND_13672(g31520,g29879,g23507);
  and AND_13673(g31523,g7528,g29333);
  and AND_13674(g31524,g29897,g20593);
  and AND_13675(g31525,g29892,g23526);
  and AND_13676(g31526,g22521,g29342);
  and AND_13677(g31527,g7553,g29343);
  and AND_13678(g31528,g19050,g29814);
  and AND_13679(g31540,g29904,g23548);
  and AND_13680(g31541,g22536,g29348);
  and AND_13681(g31542,g19050,g29814);
  and AND_13682(g31554,g19050,g29814);
  and AND_13683(g31566,g19050,g29814);
  and AND_13684(g31579,g19128,g29814);
  and AND_13685(g31654,g29325,g13062);
  and AND_13686(g31672,g29814,g19050);
  and AND_13687(g31707,g30081,g23886);
  and AND_13688(g31710,g29814,g19128);
  and AND_13689(g31744,g30092,g23902);
  and AND_13690(g31746,g30093,g23905);
  and AND_13691(g31750,g30103,g23925);
  and AND_13692(g31752,g30104,g23928);
  and AND_13693(g31756,g30114,g23942);
  and AND_13694(g31758,g30115,g23945);
  and AND_13695(g31759,g21291,g29385);
  and AND_13696(g31763,g30127,g23965);
  and AND_13697(g31765,g30128,g23968);
  and AND_13698(g31769,g30141,g23986);
  and AND_13699(g31776,g21329,g29385);
  and AND_13700(g31777,g21343,g29385);
  and AND_13701(g31778,g21369,g29385);
  and AND_13702(g31780,g30163,g23999);
  and AND_13703(g31784,g30176,g24003);
  and AND_13704(g31786,g30189,g24010);
  and AND_13705(g31787,g21281,g29385);
  and AND_13706(g31788,g21352,g29385);
  and AND_13707(g31789,g30201,g24013);
  and AND_13708(g31790,g21299,g29385);
  and AND_13709(g31792,g30214,g24017);
  and AND_13710(g31933,g939,g30735);
  and AND_13711(g31934,g31670,g18827);
  and AND_13712(g31936,g31213,g24005);
  and AND_13713(g31940,g943,g30735);
  and AND_13714(g31941,g1283,g30825);
  and AND_13715(g31943,g4717,g30614);
  and AND_13716(g31944,g31745,g22146);
  and AND_13717(g31948,g30670,g18884);
  and AND_13718(g31949,g1287,g30825);
  and AND_13719(g31959,g4907,g30673);
  and AND_13720(g31960,g31749,g22153);
  and AND_13721(g31961,g31751,g22154);
  and AND_13722(g31962,g8033,g31013);
  and AND_13723(g31963,g30731,g18895);
  and AND_13724(g31966,g31754,g22166);
  and AND_13725(g31967,g31755,g22167);
  and AND_13726(g31968,g31757,g22168);
  and AND_13727(g31969,g31189,g22139);
  and AND_13728(g31974,g31760,g22176);
  and AND_13729(g31975,g31761,g22177);
  and AND_13730(g31976,g31762,g22178);
  and AND_13731(g31977,g31764,g22179);
  and AND_13732(g31985,g4722,g30614);
  and AND_13733(g31986,g31766,g22197);
  and AND_13734(g31987,g31767,g22198);
  and AND_13735(g31988,g31768,g22199);
  and AND_13736(g31989,g31770,g22200);
  and AND_13737(g31990,g31772,g18945);
  and AND_13738(g31991,g4912,g30673);
  and AND_13739(g31992,g31773,g22213);
  and AND_13740(g31993,g31774,g22214);
  and AND_13741(g31994,g31775,g22215);
  and AND_13742(g31995,g28274,g30569);
  and AND_13743(g31996,g31779,g18979);
  and AND_13744(g32008,g31781,g22223);
  and AND_13745(g32009,g31782,g22224);
  and AND_13746(g32010,g31785,g22303);
  and AND_13747(g32011,g8287,g31134);
  and AND_13748(g32012,g8297,g31233);
  and AND_13749(g32013,g8673,g30614);
  and AND_13750(g32014,g8715,g30673);
  and AND_13751(g32016,g8522,g31138);
  and AND_13752(g32018,g4146,g30937);
  and AND_13753(g32019,g30579,g22358);
  and AND_13754(g32020,g4157,g30937);
  and AND_13755(g32028,g30569,g29339);
  and AND_13756(g32029,g31318,g16482);
  and AND_13757(g32030,g4172,g30937);
  and AND_13758(g32031,g31372,g13464);
  and AND_13759(g32032,g31373,g16515);
  and AND_13760(g32034,g14124,g31239);
  and AND_13761(g32035,g4176,g30937);
  and AND_13762(g32036,g31469,g13486);
  and AND_13763(g32039,g31476,g20070);
  and AND_13764(g32040,g14122,g31243);
  and AND_13765(g32041,g13913,g31262);
  and AND_13766(g32042,g27244,g31070);
  and AND_13767(g32043,g31482,g16173);
  and AND_13768(g32044,g31483,g20085);
  and AND_13769(g32045,g31491,g16187);
  and AND_13770(g32046,g10925,g30735);
  and AND_13771(g32047,g27248,g31070);
  and AND_13772(g32048,g31498,g13869);
  and AND_13773(g32049,g10902,g30735);
  and AND_13774(g32050,g11003,g30825);
  and AND_13775(g32051,g31506,g10831);
  and AND_13776(g32052,g31507,g13885);
  and AND_13777(g32053,g14176,g31509);
  and AND_13778(g32054,g10890,g30735);
  and AND_13779(g32055,g10999,g30825);
  and AND_13780(g32056,g27271,g31021);
  and AND_13781(g32067,g4727,g30614);
  and AND_13782(g32068,g31515,g10862);
  and AND_13783(g32069,g10878,g30735);
  and AND_13784(g32070,g10967,g30825);
  and AND_13785(g32071,g27236,g31070);
  and AND_13786(g32082,g4917,g30673);
  and AND_13787(g32083,g947,g30735);
  and AND_13788(g32084,g10948,g30825);
  and AND_13789(g32085,g27253,g31021);
  and AND_13790(g32086,g7597,g30735);
  and AND_13791(g32087,g1291,g30825);
  and AND_13792(g32088,g27241,g31070);
  and AND_13793(g32089,g27261,g31021);
  and AND_13794(g32095,g7619,g30825);
  and AND_13795(g32096,g31601,g29893);
  and AND_13796(g32097,g25960,g31021);
  and AND_13797(g32098,g4732,g30614);
  and AND_13798(g32103,g31609,g29905);
  and AND_13799(g32104,g31616,g29906);
  and AND_13800(g32105,g4922,g30673);
  and AND_13801(g32106,g31601,g29911);
  and AND_13802(g32107,g31624,g29912);
  and AND_13803(g32108,g31631,g29913);
  and AND_13804(g32109,g31609,g29920);
  and AND_13805(g32110,g31639,g29921);
  and AND_13806(g32111,g31616,g29922);
  and AND_13807(g32112,g31646,g29923);
  and AND_13808(g32113,g31601,g29925);
  and AND_13809(g32114,g31624,g29927);
  and AND_13810(g32115,g31631,g29928);
  and AND_13811(g32116,g31658,g29929);
  and AND_13812(g32119,g31609,g29939);
  and AND_13813(g32120,g31639,g29941);
  and AND_13814(g32121,g31616,g29942);
  and AND_13815(g32122,g31646,g29944);
  and AND_13816(g32126,g31601,g29948);
  and AND_13817(g32127,g31624,g29950);
  and AND_13818(g32128,g31631,g29953);
  and AND_13819(g32129,g31658,g29955);
  and AND_13820(g32139,g31601,g29960);
  and AND_13821(g32140,g31609,g29961);
  and AND_13822(g32141,g31639,g29963);
  and AND_13823(g32142,g31616,g29965);
  and AND_13824(g32143,g31646,g29967);
  and AND_13825(g32145,g31609,g29977);
  and AND_13826(g32146,g31624,g29978);
  and AND_13827(g32147,g31616,g29980);
  and AND_13828(g32148,g31631,g29981);
  and AND_13829(g32149,g31658,g29983);
  and AND_13830(g32150,g31624,g29995);
  and AND_13831(g32151,g31639,g29996);
  and AND_13832(g32152,g31631,g29998);
  and AND_13833(g32153,g31646,g29999);
  and AND_13834(g32154,g31277,g14184);
  and AND_13835(g32156,g31639,g30018);
  and AND_13836(g32157,g31646,g30021);
  and AND_13837(g32158,g31658,g30022);
  and AND_13838(g32159,g31658,g30040);
  and AND_13839(g32160,g31001,g22995);
  and AND_13840(g32161,g3151,g31154);
  and AND_13841(g32162,g31002,g23014);
  and AND_13842(g32163,g3502,g31170);
  and AND_13843(g32164,g30733,g25171);
  and AND_13844(g32165,g31669,g27742);
  and AND_13845(g32166,g31007,g23029);
  and AND_13846(g32167,g3853,g31194);
  and AND_13847(g32168,g30597,g25185);
  and AND_13848(g32169,g31014,g23046);
  and AND_13849(g32170,g31671,g27779);
  and AND_13850(g32171,g31706,g27800);
  and AND_13851(g32172,g2767,g31608);
  and AND_13852(g32173,g160,g31134);
  and AND_13853(g32174,g31708,g27837);
  and AND_13854(g32175,g31709,g27858);
  and AND_13855(g32176,g2779,g31623);
  and AND_13856(g32177,g30608,g25214);
  and AND_13857(g32178,g31747,g27886);
  and AND_13858(g32179,g31748,g27907);
  and AND_13859(g32180,g2791,g31638);
  and AND_13860(g32181,g31020,g19912);
  and AND_13861(g32182,g31753,g27937);
  and AND_13862(g32183,g2795,g31653);
  and AND_13863(g32184,g30611,g25249);
  and AND_13864(g32187,g30672,g25287);
  and AND_13865(g32188,g27586,g31376);
  and AND_13866(g32189,g30824,g25369);
  and AND_13867(g32190,g142,g31233);
  and AND_13868(g32191,g27593,g31376);
  and AND_13869(g32193,g30732,g25410);
  and AND_13870(g32194,g30601,g28436);
  and AND_13871(g32195,g30734,g25451);
  and AND_13872(g32196,g27587,g31376);
  and AND_13873(g32197,g31144,g20088);
  and AND_13874(g32198,g4253,g31327);
  and AND_13875(g32199,g30916,g25506);
  and AND_13876(g32200,g27468,g31376);
  and AND_13877(g32203,g4249,g31327);
  and AND_13878(g32204,g4245,g31327);
  and AND_13879(g32205,g30922,g28463);
  and AND_13880(g32206,g30609,g25524);
  and AND_13881(g32207,g31221,g23323);
  and AND_13882(g32224,g4300,g31327);
  and AND_13883(g32232,g31241,g20266);
  and AND_13884(g32234,g31601,g30292);
  and AND_13885(g32241,g31244,g20323);
  and AND_13886(g32242,g31245,g20324);
  and AND_13887(g32244,g31609,g30297);
  and AND_13888(g32246,g31246,g20326);
  and AND_13889(g32248,g31616,g30299);
  and AND_13890(g32254,g31247,g20379);
  and AND_13891(g32255,g31248,g20381);
  and AND_13892(g32256,g31249,g20382);
  and AND_13893(g32258,g31624,g30303);
  and AND_13894(g32260,g31250,g20385);
  and AND_13895(g32261,g31251,g20386);
  and AND_13896(g32263,g31631,g30306);
  and AND_13897(g32265,g2799,g30567);
  and AND_13898(g32269,g31253,g20443);
  and AND_13899(g32270,g31254,g20444);
  and AND_13900(g32272,g31639,g30310);
  and AND_13901(g32273,g31255,g20446);
  and AND_13902(g32274,g31256,g20447);
  and AND_13903(g32276,g31646,g30313);
  and AND_13904(g32278,g2811,g30572);
  and AND_13905(g32281,g31257,g20500);
  and AND_13906(g32282,g31258,g20503);
  and AND_13907(g32283,g31259,g20506);
  and AND_13908(g32284,g31260,g20507);
  and AND_13909(g32286,g31658,g29312);
  and AND_13910(g32287,g2823,g30578);
  and AND_13911(g32290,g31267,g20525);
  and AND_13912(g32291,g31268,g20527);
  and AND_13913(g32292,g31269,g20530);
  and AND_13914(g32293,g2827,g30593);
  and AND_13915(g32295,g27931,g31376);
  and AND_13916(g32300,g31274,g20544);
  and AND_13917(g32301,g31276,g20547);
  and AND_13918(g32302,g31279,g23485);
  and AND_13919(g32303,g27550,g31376);
  and AND_13920(g32304,g31284,g20564);
  and AND_13921(g32305,g31287,g20567);
  and AND_13922(g32306,g31289,g23499);
  and AND_13923(g32307,g31291,g23500);
  and AND_13924(g32308,g31293,g23503);
  and AND_13925(g32309,g5160,g31528);
  and AND_13926(g32310,g27577,g31376);
  and AND_13927(g32311,g31295,g20582);
  and AND_13928(g32312,g31302,g20591);
  and AND_13929(g32313,g31303,g23515);
  and AND_13930(g32314,g31304,g23516);
  and AND_13931(g32315,g31306,g23517);
  and AND_13932(g32316,g31307,g23522);
  and AND_13933(g32317,g5507,g31542);
  and AND_13934(g32321,g27613,g31376);
  and AND_13935(g32322,g31308,g20605);
  and AND_13936(g32323,g31311,g20610);
  and AND_13937(g32324,g31315,g23537);
  and AND_13938(g32325,g31316,g23538);
  and AND_13939(g32326,g31317,g23539);
  and AND_13940(g32327,g31319,g23544);
  and AND_13941(g32328,g5853,g31554);
  and AND_13942(g32330,g31320,g20631);
  and AND_13943(g32331,g31322,g20637);
  and AND_13944(g32332,g31325,g23558);
  and AND_13945(g32333,g31326,g23559);
  and AND_13946(g32334,g31375,g23568);
  and AND_13947(g32335,g6199,g31566);
  and AND_13948(g32336,g31596,g11842);
  and AND_13949(g32337,g31465,g20663);
  and AND_13950(g32338,g31466,g20668);
  and AND_13951(g32339,g31474,g20672);
  and AND_13952(g32340,g31468,g23585);
  and AND_13953(g32341,g31472,g23610);
  and AND_13954(g32342,g6545,g31579);
  and AND_13955(g32343,g31473,g20710);
  and AND_13956(g32345,g2138,g31672);
  and AND_13957(g32348,g2145,g31672);
  and AND_13958(g32350,g2697,g31710);
  and AND_13959(g32356,g2704,g31710);
  and AND_13960(g32369,g2130,g31672);
  and AND_13961(g32376,g2689,g31710);
  and AND_13962(g32396,g4698,g30983);
  and AND_13963(g32397,g31068,g15830);
  and AND_13964(g32400,g4743,g30989);
  and AND_13965(g32401,g31116,g13432);
  and AND_13966(g32402,g4888,g30990);
  and AND_13967(g32403,g31117,g15842);
  and AND_13968(g32409,g4754,g30996);
  and AND_13969(g32410,g4933,g30997);
  and AND_13970(g32411,g31119,g13469);
  and AND_13971(g32412,g4765,g30998);
  and AND_13972(g32413,g31121,g19518);
  and AND_13973(g32414,g4944,g30999);
  and AND_13974(g32418,g31126,g16239);
  and AND_13975(g32419,g4955,g31000);
  and AND_13976(g32420,g31127,g19533);
  and AND_13977(g32425,g31668,g21604);
  and AND_13978(g32428,g31133,g16261);
  and AND_13979(g33071,g31591,g32404);
  and AND_13980(g33073,g32386,g18828);
  and AND_13981(g33074,g32387,g18830);
  and AND_13982(g33081,g32388,g18875);
  and AND_13983(g33082,g32389,g18877);
  and AND_13984(g33086,g32390,g18887);
  and AND_13985(g33087,g32391,g18888);
  and AND_13986(g33091,g32392,g18897);
  and AND_13987(g33099,g32395,g18944);
  and AND_13988(g33101,g32398,g18976);
  and AND_13989(g33102,g32399,g18978);
  and AND_13990(g33104,g26296,g32137);
  and AND_13991(g33105,g26298,g32138);
  and AND_13992(g33106,g32408,g18990);
  and AND_13993(g33110,g32404,g32415);
  and AND_13994(g33111,g24005,g32421);
  and AND_13995(g33113,g31964,g22339);
  and AND_13996(g33114,g22139,g31945);
  and AND_13997(g33121,g8748,g32212);
  and AND_13998(g33122,g8859,g32192);
  and AND_13999(g33124,g8945,g32296);
  and AND_14000(g33126,g9044,g32201);
  and AND_14001(g33186,g32037,g22830);
  and AND_14002(g33233,g32094,g23005);
  and AND_14003(g33237,g32394,g25198);
  and AND_14004(g33239,g32117,g19902);
  and AND_14005(g33241,g32173,g23128);
  and AND_14006(g33242,g32123,g19931);
  and AND_14007(g33243,g32124,g19947);
  and AND_14008(g33244,g32190,g23152);
  and AND_14009(g33245,g32125,g19961);
  and AND_14010(g33247,g32130,g19980);
  and AND_14011(g33248,g32131,g19996);
  and AND_14012(g33249,g32144,g20026);
  and AND_14013(g33252,g32155,g20064);
  and AND_14014(g33263,g32393,g25481);
  and AND_14015(g33264,g31965,g21306);
  and AND_14016(g33269,g31970,g15582);
  and AND_14017(g33304,g32427,g31971);
  and AND_14018(g33305,g31935,g17811);
  and AND_14019(g33311,g31942,g12925);
  and AND_14020(g33322,g32202,g20450);
  and AND_14021(g33327,g32208,g20561);
  and AND_14022(g33328,g32209,g20584);
  and AND_14023(g33329,g32210,g20585);
  and AND_14024(g33330,g32211,g20588);
  and AND_14025(g33331,g32216,g20607);
  and AND_14026(g33332,g32217,g20608);
  and AND_14027(g33333,g32218,g20612);
  and AND_14028(g33334,g32219,g20613);
  and AND_14029(g33338,g32220,g20633);
  and AND_14030(g33339,g32221,g20634);
  and AND_14031(g33340,g32222,g20639);
  and AND_14032(g33341,g32223,g20640);
  and AND_14033(g33342,g32226,g20660);
  and AND_14034(g33343,g32227,g20665);
  and AND_14035(g33344,g32228,g20670);
  and AND_14036(g33345,g32229,g20671);
  and AND_14037(g33349,g32233,g20699);
  and AND_14038(g33350,g32235,g20702);
  and AND_14039(g33351,g32236,g20707);
  and AND_14040(g33352,g32237,g20712);
  and AND_14041(g33353,g32240,g20732);
  and AND_14042(g33355,g32243,g20769);
  and AND_14043(g33356,g32245,g20772);
  and AND_14044(g33357,g32247,g20775);
  and AND_14045(g33358,g32249,g20778);
  and AND_14046(g33359,g32252,g20853);
  and AND_14047(g33360,g32253,g20869);
  and AND_14048(g33361,g32257,g20911);
  and AND_14049(g33362,g32259,g20914);
  and AND_14050(g33363,g32262,g20918);
  and AND_14051(g33364,g32264,g20921);
  and AND_14052(g33365,g32267,g20994);
  and AND_14053(g33366,g32268,g21010);
  and AND_14054(g33367,g32271,g21053);
  and AND_14055(g33368,g32275,g21057);
  and AND_14056(g33369,g32277,g21060);
  and AND_14057(g33370,g32279,g21139);
  and AND_14058(g33371,g32280,g21155);
  and AND_14059(g33372,g32285,g21183);
  and AND_14060(g33373,g32288,g21205);
  and AND_14061(g33374,g32289,g21221);
  and AND_14062(g33376,g32294,g21268);
  and AND_14063(g33379,g30984,g32364);
  and AND_14064(g33381,g11842,g32318);
  and AND_14065(g33392,g32344,g21362);
  and AND_14066(g33399,g32346,g21379);
  and AND_14067(g33400,g32347,g21380);
  and AND_14068(g33401,g32349,g21381);
  and AND_14069(g33402,g32351,g21395);
  and AND_14070(g33403,g32352,g21396);
  and AND_14071(g33404,g32353,g21397);
  and AND_14072(g33405,g32354,g21398);
  and AND_14073(g33406,g32355,g21399);
  and AND_14074(g33407,g32357,g21406);
  and AND_14075(g33408,g32358,g21407);
  and AND_14076(g33409,g32359,g21408);
  and AND_14077(g33410,g32360,g21409);
  and AND_14078(g33411,g32361,g21410);
  and AND_14079(g33412,g32362,g21411);
  and AND_14080(g33414,g32367,g21421);
  and AND_14081(g33415,g32368,g21422);
  and AND_14082(g33416,g32370,g21423);
  and AND_14083(g33417,g32371,g21424);
  and AND_14084(g33418,g32372,g21425);
  and AND_14085(g33420,g32373,g21454);
  and AND_14086(g33421,g32374,g21455);
  and AND_14087(g33422,g32375,g21456);
  and AND_14088(g33423,g32225,g29657);
  and AND_14089(g33425,g32380,g21466);
  and AND_14090(g33428,g32230,g29672);
  and AND_14091(g33429,g32231,g29676);
  and AND_14092(g33431,g32364,g32377);
  and AND_14093(g33433,g32238,g29694);
  and AND_14094(g33434,g32239,g29702);
  and AND_14095(g33440,g32250,g29719);
  and AND_14096(g33441,g32251,g29722);
  and AND_14097(g33446,g32385,g21607);
  and AND_14098(g33450,g32266,g29737);
  and AND_14099(I31001,g29385,g32456,g32457,g32458);
  and AND_14100(I31002,g32459,g32460,g32461,g32462);
  and AND_14101(g33461,g32463,I31001,I31002);
  and AND_14102(I31006,g31376,g31796,g32464,g32465);
  and AND_14103(I31007,g32466,g32467,g32468,g32469);
  and AND_14104(g33462,g32470,I31006,I31007);
  and AND_14105(I31011,g30735,g31797,g32471,g32472);
  and AND_14106(I31012,g32473,g32474,g32475,g32476);
  and AND_14107(g33463,g32477,I31011,I31012);
  and AND_14108(I31016,g30825,g31798,g32478,g32479);
  and AND_14109(I31017,g32480,g32481,g32482,g32483);
  and AND_14110(g33464,g32484,I31016,I31017);
  and AND_14111(I31021,g31070,g31799,g32485,g32486);
  and AND_14112(I31022,g32487,g32488,g32489,g32490);
  and AND_14113(g33465,g32491,I31021,I31022);
  and AND_14114(I31026,g31194,g31800,g32492,g32493);
  and AND_14115(I31027,g32494,g32495,g32496,g32497);
  and AND_14116(g33466,g32498,I31026,I31027);
  and AND_14117(I31031,g30614,g31801,g32499,g32500);
  and AND_14118(I31032,g32501,g32502,g32503,g32504);
  and AND_14119(g33467,g32505,I31031,I31032);
  and AND_14120(I31036,g30673,g31802,g32506,g32507);
  and AND_14121(I31037,g32508,g32509,g32510,g32511);
  and AND_14122(g33468,g32512,I31036,I31037);
  and AND_14123(I31041,g31566,g31803,g32513,g32514);
  and AND_14124(I31042,g32515,g32516,g32517,g32518);
  and AND_14125(g33469,g32519,I31041,I31042);
  and AND_14126(I31046,g29385,g32521,g32522,g32523);
  and AND_14127(I31047,g32524,g32525,g32526,g32527);
  and AND_14128(g33470,g32528,I31046,I31047);
  and AND_14129(I31051,g31376,g31804,g32529,g32530);
  and AND_14130(I31052,g32531,g32532,g32533,g32534);
  and AND_14131(g33471,g32535,I31051,I31052);
  and AND_14132(I31056,g30735,g31805,g32536,g32537);
  and AND_14133(I31057,g32538,g32539,g32540,g32541);
  and AND_14134(g33472,g32542,I31056,I31057);
  and AND_14135(I31061,g30825,g31806,g32543,g32544);
  and AND_14136(I31062,g32545,g32546,g32547,g32548);
  and AND_14137(g33473,g32549,I31061,I31062);
  and AND_14138(I31066,g31070,g31807,g32550,g32551);
  and AND_14139(I31067,g32552,g32553,g32554,g32555);
  and AND_14140(g33474,g32556,I31066,I31067);
  and AND_14141(I31071,g31170,g31808,g32557,g32558);
  and AND_14142(I31072,g32559,g32560,g32561,g32562);
  and AND_14143(g33475,g32563,I31071,I31072);
  and AND_14144(I31076,g30614,g31809,g32564,g32565);
  and AND_14145(I31077,g32566,g32567,g32568,g32569);
  and AND_14146(g33476,g32570,I31076,I31077);
  and AND_14147(I31081,g30673,g31810,g32571,g32572);
  and AND_14148(I31082,g32573,g32574,g32575,g32576);
  and AND_14149(g33477,g32577,I31081,I31082);
  and AND_14150(I31086,g31554,g31811,g32578,g32579);
  and AND_14151(I31087,g32580,g32581,g32582,g32583);
  and AND_14152(g33478,g32584,I31086,I31087);
  and AND_14153(I31091,g29385,g32586,g32587,g32588);
  and AND_14154(I31092,g32589,g32590,g32591,g32592);
  and AND_14155(g33479,g32593,I31091,I31092);
  and AND_14156(I31096,g31376,g31812,g32594,g32595);
  and AND_14157(I31097,g32596,g32597,g32598,g32599);
  and AND_14158(g33480,g32600,I31096,I31097);
  and AND_14159(I31101,g30735,g31813,g32601,g32602);
  and AND_14160(I31102,g32603,g32604,g32605,g32606);
  and AND_14161(g33481,g32607,I31101,I31102);
  and AND_14162(I31106,g30825,g31814,g32608,g32609);
  and AND_14163(I31107,g32610,g32611,g32612,g32613);
  and AND_14164(g33482,g32614,I31106,I31107);
  and AND_14165(I31111,g31070,g31815,g32615,g32616);
  and AND_14166(I31112,g32617,g32618,g32619,g32620);
  and AND_14167(g33483,g32621,I31111,I31112);
  and AND_14168(I31116,g31154,g31816,g32622,g32623);
  and AND_14169(I31117,g32624,g32625,g32626,g32627);
  and AND_14170(g33484,g32628,I31116,I31117);
  and AND_14171(I31121,g30614,g31817,g32629,g32630);
  and AND_14172(I31122,g32631,g32632,g32633,g32634);
  and AND_14173(g33485,g32635,I31121,I31122);
  and AND_14174(I31126,g30673,g31818,g32636,g32637);
  and AND_14175(I31127,g32638,g32639,g32640,g32641);
  and AND_14176(g33486,g32642,I31126,I31127);
  and AND_14177(I31131,g31542,g31819,g32643,g32644);
  and AND_14178(I31132,g32645,g32646,g32647,g32648);
  and AND_14179(g33487,g32649,I31131,I31132);
  and AND_14180(I31136,g29385,g32651,g32652,g32653);
  and AND_14181(I31137,g32654,g32655,g32656,g32657);
  and AND_14182(g33488,g32658,I31136,I31137);
  and AND_14183(I31141,g31376,g31820,g32659,g32660);
  and AND_14184(I31142,g32661,g32662,g32663,g32664);
  and AND_14185(g33489,g32665,I31141,I31142);
  and AND_14186(I31146,g30735,g31821,g32666,g32667);
  and AND_14187(I31147,g32668,g32669,g32670,g32671);
  and AND_14188(g33490,g32672,I31146,I31147);
  and AND_14189(I31151,g30825,g31822,g32673,g32674);
  and AND_14190(I31152,g32675,g32676,g32677,g32678);
  and AND_14191(g33491,g32679,I31151,I31152);
  and AND_14192(I31156,g31070,g31823,g32680,g32681);
  and AND_14193(I31157,g32682,g32683,g32684,g32685);
  and AND_14194(g33492,g32686,I31156,I31157);
  and AND_14195(I31161,g30614,g31824,g32687,g32688);
  and AND_14196(I31162,g32689,g32690,g32691,g32692);
  and AND_14197(g33493,g32693,I31161,I31162);
  and AND_14198(I31166,g30673,g31825,g32694,g32695);
  and AND_14199(I31167,g32696,g32697,g32698,g32699);
  and AND_14200(g33494,g32700,I31166,I31167);
  and AND_14201(I31171,g31528,g31826,g32701,g32702);
  and AND_14202(I31172,g32703,g32704,g32705,g32706);
  and AND_14203(g33495,g32707,I31171,I31172);
  and AND_14204(I31176,g31579,g31827,g32708,g32709);
  and AND_14205(I31177,g32710,g32711,g32712,g32713);
  and AND_14206(g33496,g32714,I31176,I31177);
  and AND_14207(I31181,g29385,g32716,g32717,g32718);
  and AND_14208(I31182,g32719,g32720,g32721,g32722);
  and AND_14209(g33497,g32723,I31181,I31182);
  and AND_14210(I31186,g31376,g31828,g32724,g32725);
  and AND_14211(I31187,g32726,g32727,g32728,g32729);
  and AND_14212(g33498,g32730,I31186,I31187);
  and AND_14213(I31191,g30735,g31829,g32731,g32732);
  and AND_14214(I31192,g32733,g32734,g32735,g32736);
  and AND_14215(g33499,g32737,I31191,I31192);
  and AND_14216(I31196,g30825,g31830,g32738,g32739);
  and AND_14217(I31197,g32740,g32741,g32742,g32743);
  and AND_14218(g33500,g32744,I31196,I31197);
  and AND_14219(I31201,g31672,g31831,g32745,g32746);
  and AND_14220(I31202,g32747,g32748,g32749,g32750);
  and AND_14221(g33501,g32751,I31201,I31202);
  and AND_14222(I31206,g31710,g31832,g32752,g32753);
  and AND_14223(I31207,g32754,g32755,g32756,g32757);
  and AND_14224(g33502,g32758,I31206,I31207);
  and AND_14225(I31211,g31021,g31833,g32759,g32760);
  and AND_14226(I31212,g32761,g32762,g32763,g32764);
  and AND_14227(g33503,g32765,I31211,I31212);
  and AND_14228(I31216,g30937,g31834,g32766,g32767);
  and AND_14229(I31217,g32768,g32769,g32770,g32771);
  and AND_14230(g33504,g32772,I31216,I31217);
  and AND_14231(I31221,g31327,g31835,g32773,g32774);
  and AND_14232(I31222,g32775,g32776,g32777,g32778);
  and AND_14233(g33505,g32779,I31221,I31222);
  and AND_14234(I31226,g29385,g32781,g32782,g32783);
  and AND_14235(I31227,g32784,g32785,g32786,g32787);
  and AND_14236(g33506,g32788,I31226,I31227);
  and AND_14237(I31231,g31376,g31836,g32789,g32790);
  and AND_14238(I31232,g32791,g32792,g32793,g32794);
  and AND_14239(g33507,g32795,I31231,I31232);
  and AND_14240(I31236,g30735,g31837,g32796,g32797);
  and AND_14241(I31237,g32798,g32799,g32800,g32801);
  and AND_14242(g33508,g32802,I31236,I31237);
  and AND_14243(I31241,g30825,g31838,g32803,g32804);
  and AND_14244(I31242,g32805,g32806,g32807,g32808);
  and AND_14245(g33509,g32809,I31241,I31242);
  and AND_14246(I31246,g31672,g31839,g32810,g32811);
  and AND_14247(I31247,g32812,g32813,g32814,g32815);
  and AND_14248(g33510,g32816,I31246,I31247);
  and AND_14249(I31251,g31710,g31840,g32817,g32818);
  and AND_14250(I31252,g32819,g32820,g32821,g32822);
  and AND_14251(g33511,g32823,I31251,I31252);
  and AND_14252(I31256,g31021,g31841,g32824,g32825);
  and AND_14253(I31257,g32826,g32827,g32828,g32829);
  and AND_14254(g33512,g32830,I31256,I31257);
  and AND_14255(I31261,g30937,g31842,g32831,g32832);
  and AND_14256(I31262,g32833,g32834,g32835,g32836);
  and AND_14257(g33513,g32837,I31261,I31262);
  and AND_14258(I31266,g31327,g31843,g32838,g32839);
  and AND_14259(I31267,g32840,g32841,g32842,g32843);
  and AND_14260(g33514,g32844,I31266,I31267);
  and AND_14261(I31271,g29385,g32846,g32847,g32848);
  and AND_14262(I31272,g32849,g32850,g32851,g32852);
  and AND_14263(g33515,g32853,I31271,I31272);
  and AND_14264(I31276,g31376,g31844,g32854,g32855);
  and AND_14265(I31277,g32856,g32857,g32858,g32859);
  and AND_14266(g33516,g32860,I31276,I31277);
  and AND_14267(I31281,g30735,g31845,g32861,g32862);
  and AND_14268(I31282,g32863,g32864,g32865,g32866);
  and AND_14269(g33517,g32867,I31281,I31282);
  and AND_14270(I31286,g30825,g31846,g32868,g32869);
  and AND_14271(I31287,g32870,g32871,g32872,g32873);
  and AND_14272(g33518,g32874,I31286,I31287);
  and AND_14273(I31291,g31021,g31847,g32875,g32876);
  and AND_14274(I31292,g32877,g32878,g32879,g32880);
  and AND_14275(g33519,g32881,I31291,I31292);
  and AND_14276(I31296,g30937,g31848,g32882,g32883);
  and AND_14277(I31297,g32884,g32885,g32886,g32887);
  and AND_14278(g33520,g32888,I31296,I31297);
  and AND_14279(I31301,g31327,g31849,g32889,g32890);
  and AND_14280(I31302,g32891,g32892,g32893,g32894);
  and AND_14281(g33521,g32895,I31301,I31302);
  and AND_14282(I31306,g30614,g31850,g32896,g32897);
  and AND_14283(I31307,g32898,g32899,g32900,g32901);
  and AND_14284(g33522,g32902,I31306,I31307);
  and AND_14285(I31311,g30673,g31851,g32903,g32904);
  and AND_14286(I31312,g32905,g32906,g32907,g32908);
  and AND_14287(g33523,g32909,I31311,I31312);
  and AND_14288(I31316,g29385,g32911,g32912,g32913);
  and AND_14289(I31317,g32914,g32915,g32916,g32917);
  and AND_14290(g33524,g32918,I31316,I31317);
  and AND_14291(I31321,g31376,g31852,g32919,g32920);
  and AND_14292(I31322,g32921,g32922,g32923,g32924);
  and AND_14293(g33525,g32925,I31321,I31322);
  and AND_14294(I31326,g30735,g31853,g32926,g32927);
  and AND_14295(I31327,g32928,g32929,g32930,g32931);
  and AND_14296(g33526,g32932,I31326,I31327);
  and AND_14297(I31331,g30825,g31854,g32933,g32934);
  and AND_14298(I31332,g32935,g32936,g32937,g32938);
  and AND_14299(g33527,g32939,I31331,I31332);
  and AND_14300(I31336,g31672,g31855,g32940,g32941);
  and AND_14301(I31337,g32942,g32943,g32944,g32945);
  and AND_14302(g33528,g32946,I31336,I31337);
  and AND_14303(I31341,g31710,g31856,g32947,g32948);
  and AND_14304(I31342,g32949,g32950,g32951,g32952);
  and AND_14305(g33529,g32953,I31341,I31342);
  and AND_14306(I31346,g31021,g31857,g32954,g32955);
  and AND_14307(I31347,g32956,g32957,g32958,g32959);
  and AND_14308(g33530,g32960,I31346,I31347);
  and AND_14309(I31351,g30937,g31858,g32961,g32962);
  and AND_14310(I31352,g32963,g32964,g32965,g32966);
  and AND_14311(g33531,g32967,I31351,I31352);
  and AND_14312(I31356,g31327,g31859,g32968,g32969);
  and AND_14313(I31357,g32970,g32971,g32972,g32973);
  and AND_14314(g33532,g32974,I31356,I31357);
  and AND_14315(g33639,g33386,g18829);
  and AND_14316(g33640,g33387,g18831);
  and AND_14317(g33646,g33389,g18876);
  and AND_14318(g33647,g33390,g18878);
  and AND_14319(g33652,g33393,g18889);
  and AND_14320(g33657,g30991,g33443);
  and AND_14321(g33674,g33164,g10710,g22319);
  and AND_14322(g33675,g33164,g10727,g22332);
  and AND_14323(g33676,g33125,g7970);
  and AND_14324(g33677,g33443,g31937);
  and AND_14325(g33678,g33149,g10710,g22319);
  and AND_14326(g33680,g33128,g4688);
  and AND_14327(g33681,g33129,g7991);
  and AND_14328(g33683,g33149,g10727,g22332);
  and AND_14329(g33684,g33139,g13565);
  and AND_14330(g33687,g33132,g4878);
  and AND_14331(g33689,g33144,g11006);
  and AND_14332(g33690,g33146,g16280);
  and AND_14333(g33693,g33145,g13594);
  and AND_14334(g33697,g33160,g13330);
  and AND_14335(g33700,g33148,g11012);
  and AND_14336(g33701,g33162,g16305);
  and AND_14337(g33704,g33176,g10710,g22319);
  and AND_14338(g33707,g33174,g13346);
  and AND_14339(g33710,g14037,g33246);
  and AND_14340(g33711,g33176,g10727,g22332);
  and AND_14341(g33715,g33135,g19416);
  and AND_14342(g33717,g14092,g33306);
  and AND_14343(g33718,g33147,g19432);
  and AND_14344(g33719,g33141,g19433);
  and AND_14345(g33720,g33161,g19439);
  and AND_14346(g33721,g33163,g19440);
  and AND_14347(g33722,g33175,g19445);
  and AND_14348(g33723,g14091,g33299);
  and AND_14349(g33724,g14145,g33258);
  and AND_14350(g33725,g22626,g10851,g33176);
  and AND_14351(g33727,g33115,g19499);
  and AND_14352(g33728,g22626,g10851,g33187);
  and AND_14353(g33730,g7202,g4621,g33127,g4633);
  and AND_14354(g33731,g33116,g19520);
  and AND_14355(I31593,g31003,g8350,g7788);
  and AND_14356(g33734,g7806,g33136,I31593);
  and AND_14357(g33735,g33118,g19553);
  and AND_14358(I31600,g31009,g8400,g7809);
  and AND_14359(g33742,g7828,g33142,I31600);
  and AND_14360(g33743,g33119,g19574);
  and AND_14361(g33758,g33133,g20269);
  and AND_14362(g33759,g33123,g22847);
  and AND_14363(g33760,g33143,g20328);
  and AND_14364(g33784,g33107,g20531);
  and AND_14365(g33785,g33100,g20550);
  and AND_14366(g33786,g33130,g20572);
  and AND_14367(g33787,g33103,g20595);
  and AND_14368(g33789,g33159,g23022);
  and AND_14369(g33790,g33108,g20643);
  and AND_14370(g33795,g33138,g20782);
  and AND_14371(g33796,g33117,g25267);
  and AND_14372(g33798,g33227,g20058);
  and AND_14373(g33801,g33437,g25327);
  and AND_14374(g33802,g33097,g14545);
  and AND_14375(g33803,g33231,g20071);
  and AND_14376(g33805,g33232,g20079);
  and AND_14377(g33807,g33112,g25452);
  and AND_14378(g33808,g33109,g22161);
  and AND_14379(g33809,g33432,g30184);
  and AND_14380(g33810,g33427,g12768);
  and AND_14381(g33811,g33439,g17573);
  and AND_14382(g33812,g23088,g33187,g9104);
  and AND_14383(g33814,g33098,g28144);
  and AND_14384(g33815,g33449,g12911);
  and AND_14385(g33816,g33234,g20096);
  and AND_14386(g33817,g33235,g20102);
  and AND_14387(g33818,g33236,g20113);
  and AND_14388(g33819,g23088,g33176,g9104);
  and AND_14389(g33820,g33075,g26830);
  and AND_14390(g33821,g33238,g20153);
  and AND_14391(g33822,g33385,g20157);
  and AND_14392(g33828,g33090,g24411);
  and AND_14393(g33829,g33240,g20164);
  and AND_14394(g33830,g33382,g20166);
  and AND_14395(g33831,g23088,g33149,g9104);
  and AND_14396(g33832,g33088,g27991);
  and AND_14397(g33833,g33093,g25852);
  and AND_14398(g33834,g33095,g29172);
  and AND_14399(g33835,g4340,g33413);
  and AND_14400(g33836,g33096,g27020);
  and AND_14401(g33837,g33251,g20233);
  and AND_14402(g33840,g33253,g20267);
  and AND_14403(g33841,g33254,g20268);
  and AND_14404(g33842,g33255,g20322);
  and AND_14405(g33843,g33256,g20325);
  and AND_14406(g33844,g33257,g20327);
  and AND_14407(g33846,g33259,g20380);
  and AND_14408(g33847,g33260,g20383);
  and AND_14409(g33848,g33261,g20384);
  and AND_14410(g33849,g33262,g20387);
  and AND_14411(g33855,g33265,g20441);
  and AND_14412(g33856,g33266,g20442);
  and AND_14413(g33857,g33267,g20445);
  and AND_14414(g33858,g33268,g20448);
  and AND_14415(g33859,g33426,g10531);
  and AND_14416(g33860,g33270,g20501);
  and AND_14417(g33861,g33271,g20502);
  and AND_14418(g33862,g33272,g20504);
  and AND_14419(g33863,g33273,g20505);
  and AND_14420(g33864,g33274,g20524);
  and AND_14421(g33865,g33275,g20526);
  and AND_14422(g33866,g33276,g20528);
  and AND_14423(g33867,g33277,g20529);
  and AND_14424(g33868,g33278,g20542);
  and AND_14425(g33869,g33279,g20543);
  and AND_14426(g33870,g33280,g20545);
  and AND_14427(g33871,g33281,g20546);
  and AND_14428(g33872,g33282,g20548);
  and AND_14429(g33873,g33291,g20549);
  and AND_14430(g33876,g33286,g20562);
  and AND_14431(g33877,g33287,g20563);
  and AND_14432(g33878,g33288,g20565);
  and AND_14433(g33879,g33289,g20566);
  and AND_14434(g33880,g33290,g20568);
  and AND_14435(g33881,g33292,g20586);
  and AND_14436(g33882,g33293,g20587);
  and AND_14437(g33883,g33294,g20589);
  and AND_14438(g33884,g33295,g20590);
  and AND_14439(g33885,g33296,g20609);
  and AND_14440(g33886,g33297,g20614);
  and AND_14441(g33887,g33298,g20615);
  and AND_14442(g33889,g33303,g20641);
  and AND_14443(g33890,g33310,g20659);
  and AND_14444(g33892,g33312,g20701);
  and AND_14445(g33893,g33313,g20706);
  and AND_14446(g33896,g33314,g20771);
  and AND_14447(g33897,g33315,g20777);
  and AND_14448(g33898,g33419,g15655);
  and AND_14449(g33899,g32132,g33335);
  and AND_14450(g33900,g33316,g20913);
  and AND_14451(g33901,g33317,g20920);
  and AND_14452(g33902,g33085,g13202);
  and AND_14453(g33903,g33447,g19146);
  and AND_14454(g33904,g33321,g21059);
  and AND_14455(g33905,g33089,g15574);
  and AND_14456(g33906,g33084,g22311);
  and AND_14457(g33907,g23088,g33219,g9104);
  and AND_14458(g33908,g33092,g18935);
  and AND_14459(g33909,g33131,g10708);
  and AND_14460(g33910,g33134,g7836);
  and AND_14461(g33911,g33137,g10725);
  and AND_14462(g33913,g23088,g33204,g9104);
  and AND_14463(g33915,g33140,g7846);
  and AND_14464(g33919,g33438,g10795);
  and AND_14465(g33921,g33187,g9104,g19200);
  and AND_14466(g33922,g33448,g7202);
  and AND_14467(g33924,g33335,g33346);
  and AND_14468(g33927,g33094,g21412);
  and AND_14469(g33941,g33380,g21560);
  and AND_14470(g33942,g33383,g21608);
  and AND_14471(g33943,g33384,g21609);
  and AND_14472(g34045,g33766,g22942);
  and AND_14473(g34050,g33772,g22942);
  and AND_14474(g34054,g33778,g22942);
  and AND_14475(g34061,g33800,g23076);
  and AND_14476(g34063,g33806,g23121);
  and AND_14477(g34065,g33813,g23148);
  and AND_14478(g34066,g33730,g19352);
  and AND_14479(g34069,g8774,g33797);
  and AND_14480(g34071,g8854,g33799);
  and AND_14481(g34072,g33839,g24872);
  and AND_14482(g34073,g8948,g33823);
  and AND_14483(g34074,g33685,g19498);
  and AND_14484(g34075,g33692,g19517);
  and AND_14485(g34076,g33694,g19519);
  and AND_14486(g34077,g22957,g9104,g33736);
  and AND_14487(g34078,g33699,g19531);
  and AND_14488(g34079,g33703,g19532);
  and AND_14489(g34080,g22957,g9104,g33750);
  and AND_14490(g34081,g33706,g19552);
  and AND_14491(g34082,g33709,g19554);
  and AND_14492(g34083,g33714,g19573);
  and AND_14493(g34084,g9214,g33851);
  and AND_14494(g34085,g33761,g9104,g18957);
  and AND_14495(g34086,g20114,g33766,g9104);
  and AND_14496(g34087,g33766,g9104,g18957);
  and AND_14497(g34088,g33736,g9104,g18957);
  and AND_14498(g34089,g22957,g9104,g33744);
  and AND_14499(g34091,g22957,g9104,g33761);
  and AND_14500(g34092,g33750,g9104,g18957);
  and AND_14501(g34093,g20114,g33755,g9104);
  and AND_14502(g34096,g22957,g9104,g33772);
  and AND_14503(g34097,g33772,g9104,g18957);
  and AND_14504(g34098,g33744,g9104,g18957);
  and AND_14505(g34102,g33912,g23599);
  and AND_14506(g34104,g33916,g23639);
  and AND_14507(g34105,g33778,g9104,g18957);
  and AND_14508(g34106,g33917,g23675);
  and AND_14509(g34108,g22957,g9104,g33766);
  and AND_14510(g34109,g33918,g23708);
  and AND_14511(g34110,g33732,g22935);
  and AND_14512(g34111,g33733,g22936);
  and AND_14513(g34112,g22957,g9104,g33778);
  and AND_14514(g34113,g33734,g19744);
  and AND_14515(g34114,g33920,g23742);
  and AND_14516(g34115,g20516,g9104,g33750);
  and AND_14517(g34116,g33933,g25140);
  and AND_14518(g34117,g33742,g19755);
  and AND_14519(g34119,g20516,g9104,g33755);
  and AND_14520(g34120,g33930,g25158);
  and AND_14521(g34133,g33845,g23958);
  and AND_14522(g34135,g33926,g23802);
  and AND_14523(g34136,g33850,g23293);
  and AND_14524(g34137,g33928,g23802);
  and AND_14525(g34138,g33929,g23828);
  and AND_14526(g34139,g33827,g23314);
  and AND_14527(g34140,g33931,g23802);
  and AND_14528(g34141,g33932,g23828);
  and AND_14529(g34143,g33934,g23828);
  and AND_14530(g34146,g33788,g20091);
  and AND_14531(g34157,g33794,g20159);
  and AND_14532(g34169,g33804,g31227);
  and AND_14533(g34171,g33925,g24360);
  and AND_14534(g34173,g33679,g24368);
  and AND_14535(g34178,g33712,g24361);
  and AND_14536(g34179,g33686,g24372);
  and AND_14537(g34180,g33716,g24373);
  and AND_14538(g34182,g33691,g24384);
  and AND_14539(g34183,g33695,g24385);
  and AND_14540(g34184,g33698,g24388);
  and AND_14541(g34185,g33702,g24389);
  and AND_14542(g34186,g33705,g24396);
  and AND_14543(g34187,g33708,g24397);
  and AND_14544(g34191,g33713,g24404);
  and AND_14545(g34196,g33682,g24485);
  and AND_14546(g34198,g33688,g24491);
  and AND_14547(g34203,g33726,g24537);
  and AND_14548(g34205,g33729,g24541);
  and AND_14549(g34211,g33891,g21349);
  and AND_14550(g34212,g33761,g22689);
  and AND_14551(g34213,g33766,g22689);
  and AND_14552(g34214,g33772,g22689);
  and AND_14553(g34215,g33778,g22670);
  and AND_14554(g34216,g33778,g22689);
  and AND_14555(g34217,g33736,g22876);
  and AND_14556(g34218,g33744,g22670);
  and AND_14557(g34219,g33736,g22942);
  and AND_14558(g34223,g33744,g22876);
  and AND_14559(g34224,g33736,g22670);
  and AND_14560(g34225,g33744,g22942);
  and AND_14561(g34226,g33914,g21467);
  and AND_14562(g34228,g33750,g22942);
  and AND_14563(g34230,g33761,g22942);
  and AND_14564(g34279,g34231,g19208);
  and AND_14565(g34281,g34043,g19276);
  and AND_14566(g34284,g34046,g19351);
  and AND_14567(g34287,g11370,g34124);
  and AND_14568(g34291,g34055,g19366);
  and AND_14569(g34295,g34057,g19370);
  and AND_14570(g34298,g8679,g34132);
  and AND_14571(g34301,g34064,g19415);
  and AND_14572(g34309,g13947,g34147);
  and AND_14573(g34310,g14003,g34162);
  and AND_14574(g34319,g9535,g34156);
  and AND_14575(g34322,g14188,g34174);
  and AND_14576(g34324,g14064,g34161);
  and AND_14577(g34329,g14511,g34181);
  and AND_14578(g34333,g9984,g34192);
  and AND_14579(g34334,g34090,g19865);
  and AND_14580(g34335,g8461,g34197);
  and AND_14581(g34337,g34095,g19881);
  and AND_14582(g34338,g34099,g19905);
  and AND_14583(g34340,g34100,g19950);
  and AND_14584(g34341,g34101,g19952);
  and AND_14585(g34342,g34103,g19998);
  and AND_14586(g34344,g34107,g20038);
  and AND_14587(g34348,g34125,g20128);
  and AND_14588(g34363,g34148,g20389);
  and AND_14589(g34364,g34048,g24366);
  and AND_14590(g34365,g34149,g20451);
  and AND_14591(g34367,g7404,g34042);
  and AND_14592(g34370,g34067,g10554);
  and AND_14593(g34371,g7450,g34044);
  and AND_14594(g34375,g13077,g34049);
  and AND_14595(g34378,g13095,g34053);
  and AND_14596(g34380,g34158,g20571);
  and AND_14597(g34381,g34166,g20594);
  and AND_14598(g34382,g34167,g20618);
  and AND_14599(g34385,g34168,g20642);
  and AND_14600(g34386,g10800,g34060);
  and AND_14601(g34388,g10802,g34062);
  and AND_14602(g34389,g34170,g20715);
  and AND_14603(g34390,g34172,g21069);
  and AND_14604(g34393,g34189,g21304);
  and AND_14605(g34394,g34190,g21305);
  and AND_14606(g34395,g34193,g21336);
  and AND_14607(g34396,g34194,g21337);
  and AND_14608(g34397,g7673,g34068);
  and AND_14609(g34398,g7684,g34070);
  and AND_14610(g34401,g34199,g21383);
  and AND_14611(g34410,g34204,g21427);
  and AND_14612(g34413,g34094,g22670);
  and AND_14613(g34414,g34206,g21457);
  and AND_14614(g34415,g34207,g21458);
  and AND_14615(g34470,g7834,g34325);
  and AND_14616(g34474,g20083,g34326);
  and AND_14617(g34475,g27450,g34327);
  and AND_14618(g34476,g34399,g18891);
  and AND_14619(g34477,g26344,g34328);
  and AND_14620(g34478,g34402,g18904);
  and AND_14621(g34479,g34403,g18905);
  and AND_14622(g34481,g34404,g18916);
  and AND_14623(g34482,g34405,g18917);
  and AND_14624(g34483,g34406,g18938);
  and AND_14625(g34484,g34407,g18939);
  and AND_14626(g34485,g34411,g18952);
  and AND_14627(g34486,g34412,g18953);
  and AND_14628(g34487,g34416,g18983);
  and AND_14629(g34488,g34417,g18988);
  and AND_14630(g34489,g34421,g19068);
  and AND_14631(g34492,g34272,g33430);
  and AND_14632(g34493,g34273,g19360);
  and AND_14633(g34495,g34274,g19365);
  and AND_14634(g34497,g34275,g33072);
  and AND_14635(g34498,g13888,g34336);
  and AND_14636(g34499,g31288,g34339);
  and AND_14637(g34500,g34276,g30568);
  and AND_14638(g34502,g26363,g34343);
  and AND_14639(g34503,g34278,g19437);
  and AND_14640(g34506,g8833,g34354);
  and AND_14641(g34507,g34280,g19454);
  and AND_14642(g34508,g34282,g19472);
  and AND_14643(g34509,g34283,g19473);
  and AND_14644(g34513,g9003,g34346);
  and AND_14645(g34514,g34286,g19480);
  and AND_14646(g34515,g34288,g19491);
  and AND_14647(g34516,g34289,g19492);
  and AND_14648(g34517,g34290,g19493);
  and AND_14649(g34518,g34292,g19503);
  and AND_14650(g34519,g34293,g19504);
  and AND_14651(g34520,g34294,g19505);
  and AND_14652(g34523,g9162,g34351);
  and AND_14653(g34524,g9083,g34359);
  and AND_14654(g34525,g34297,g19528);
  and AND_14655(g34526,g34300,g19569);
  and AND_14656(g34527,g34303,g19603);
  and AND_14657(g34528,g34305,g19617);
  and AND_14658(g34529,g34306,g19634);
  and AND_14659(g34532,g34314,g19710);
  and AND_14660(g34533,g34318,g19731);
  and AND_14661(g34534,g34321,g19743);
  and AND_14662(g34538,g34330,g20054);
  and AND_14663(g34541,g34331,g20087);
  and AND_14664(g34542,g34332,g20089);
  and AND_14665(g34554,g34347,g20495);
  and AND_14666(g34555,g34349,g20512);
  and AND_14667(g34556,g34350,g20537);
  and AND_14668(g34557,g34352,g20555);
  and AND_14669(g34558,g34353,g20578);
  and AND_14670(g34560,g34366,g17366);
  and AND_14671(g34561,g34368,g17410);
  and AND_14672(g34562,g34369,g17411);
  and AND_14673(g34563,g34372,g17465);
  and AND_14674(g34564,g34373,g17466);
  and AND_14675(g34565,g34374,g17471);
  and AND_14676(g34566,g34376,g17489);
  and AND_14677(g34567,g34377,g17491);
  and AND_14678(g34568,g34379,g17512);
  and AND_14679(g34571,g27225,g34299);
  and AND_14680(g34572,g34387,g33326);
  and AND_14681(g34577,g24577,g34307);
  and AND_14682(g34578,g24578,g34308);
  and AND_14683(g34580,g29539,g34311);
  and AND_14684(g34581,g22864,g34312);
  and AND_14685(g34582,g7764,g34313);
  and AND_14686(g34584,g24653,g34315);
  and AND_14687(g34585,g24705,g34316);
  and AND_14688(g34586,g11025,g34317);
  and AND_14689(g34588,g26082,g34323);
  and AND_14690(g34655,g34573,g18885);
  and AND_14691(g34658,g34574,g18896);
  and AND_14692(g34661,g34575,g18907);
  and AND_14693(g34662,g34576,g18931);
  and AND_14694(g34665,g34583,g19067);
  and AND_14695(g34666,g34587,g19144);
  and AND_14696(g34667,g34471,g33424);
  and AND_14697(g34678,g34490,g19431);
  and AND_14698(g34679,g14093,g34539);
  and AND_14699(g34681,g34491,g19438);
  and AND_14700(g34684,g14178,g34545);
  and AND_14701(g34685,g14164,g34550);
  and AND_14702(g34686,g34494,g19494);
  and AND_14703(g34687,g14181,g34543);
  and AND_14704(g34694,g34530,g19885);
  and AND_14705(g34696,g34531,g20004);
  and AND_14706(g34700,g34535,g20129);
  and AND_14707(g34701,g34536,g20179);
  and AND_14708(g34702,g34537,g20208);
  and AND_14709(g34706,g34496,g10570);
  and AND_14710(g34707,g34544,g20579);
  and AND_14711(g34709,g34549,g17242);
  and AND_14712(g34710,g34553,g20903);
  and AND_14713(g34715,g34570,g33375);
  and AND_14714(g34738,g34660,g33442);
  and AND_14715(g34740,g34664,g19414);
  and AND_14716(g34741,g8899,g34697);
  and AND_14717(g34742,g9000,g34698);
  and AND_14718(g34743,g8951,g34703);
  and AND_14719(g34744,g34668,g19481);
  and AND_14720(g34745,g34669,g19482);
  and AND_14721(g34746,g34670,g19526);
  and AND_14722(g34747,g34671,g19527);
  and AND_14723(g34748,g34672,g19529);
  and AND_14724(g34750,g34673,g19542);
  and AND_14725(g34751,g34674,g19543);
  and AND_14726(g34752,g34675,g19544);
  and AND_14727(g34753,g34676,g19586);
  and AND_14728(g34754,g34677,g19602);
  and AND_14729(g34756,g34680,g19618);
  and AND_14730(g34757,g34682,g19635);
  and AND_14731(g34758,g34683,g19657);
  and AND_14732(g34763,g34689,g19915);
  and AND_14733(g34764,g34691,g20009);
  and AND_14734(g34765,g34692,g20057);
  and AND_14735(g34771,g34693,g20147);
  and AND_14736(g34774,g34695,g20180);
  and AND_14737(g34782,g34711,g33888);
  and AND_14738(g34811,g14165,g34766);
  and AND_14739(g34841,g34761,g20080);
  and AND_14740(g34842,g34762,g20168);
  and AND_14741(g34857,g16540,g34813);
  and AND_14742(g34858,g16540,g34816);
  and AND_14743(g34859,g16540,g34820);
  and AND_14744(g34860,g16540,g34823);
  and AND_14745(g34861,g16540,g34827);
  and AND_14746(g34862,g16540,g34830);
  and AND_14747(g34863,g16540,g34833);
  and AND_14748(g34865,g16540,g34836);
  and AND_14749(g34866,g34819,g20106);
  and AND_14750(g34867,g34826,g20145);
  and AND_14751(g34868,g34813,g19866);
  and AND_14752(g34869,g34816,g19869);
  and AND_14753(g34870,g34820,g19882);
  and AND_14754(g34871,g34823,g19908);
  and AND_14755(g34872,g34827,g19954);
  and AND_14756(g34873,g34830,g20046);
  and AND_14757(g34874,g34833,g20060);
  and AND_14758(g34875,g34836,g20073);
  and AND_14759(g34876,g34844,g20534);
  and AND_14760(g34909,g34856,g20130);
  and AND_14761(g34948,g16540,g34935);
  and AND_14762(g34953,g34935,g19957);
  and AND_14763(g34955,g34931,g34320);
  and AND_14764(g34961,g34944,g23019);
  and AND_14765(g34962,g34945,g23020);
  and AND_14766(g34963,g34946,g23041);
  and AND_14767(g34964,g34947,g23060);
  and AND_14768(g34965,g34949,g23084);
  and AND_14769(g34966,g34950,g23170);
  and AND_14770(g34967,g34951,g23189);
  and AND_14771(g34968,g34952,g23203);
  and AND_14772(g34969,g34960,g19570);
  and AND_14773(g34999,g34998,g23085);
  or OR_14774(g7404,g933,g939);
  or OR_14775(g7450,g1277,g1283);
  or OR_14776(g7673,g4153,g4172);
  or OR_14777(g7684,g4072,g4176);
  or OR_14778(g7764,g2999,g2932);
  or OR_14779(g7834,g2886,g2946);
  or OR_14780(g7932,g4072,g4153);
  or OR_14781(I12583,g1157,g1239,g990);
  or OR_14782(g8417,g1056,g1116,I12583);
  or OR_14783(g8461,g301,g534);
  or OR_14784(I12611,g1500,g1582,g1333);
  or OR_14785(g8476,g1399,g1459,I12611);
  or OR_14786(g8679,g222,g199);
  or OR_14787(I12782,g4188,g4194,g4197,g4200);
  or OR_14788(I12783,g4204,g4207,g4210,g4180);
  or OR_14789(g8790,I12782,I12783);
  or OR_14790(g8863,g1644,g1664);
  or OR_14791(g8904,g1779,g1798);
  or OR_14792(g8905,g2204,g2223);
  or OR_14793(I12902,g4235,g4232,g4229,g4226);
  or OR_14794(I12903,g4222,g4219,g4216,g4213);
  or OR_14795(g8921,I12902,I12903);
  or OR_14796(g8956,g1913,g1932);
  or OR_14797(g8957,g2338,g2357);
  or OR_14798(g9012,g2047,g2066);
  or OR_14799(g9013,g2472,g2491);
  or OR_14800(g9055,g2606,g2625);
  or OR_14801(g9483,g1008,g969);
  or OR_14802(g9535,g209,g538);
  or OR_14803(g9536,g1351,g1312);
  or OR_14804(g9984,g4300,g4242);
  or OR_14805(g10589,g7223,g7201);
  or OR_14806(g10800,g7517,g952);
  or OR_14807(g10802,g7533,g1296);
  or OR_14808(g11025,g2980,g7831);
  or OR_14809(g11370,g8807,g550);
  or OR_14810(g11372,g490,g482,g8038);
  or OR_14811(g11380,g8583,g8530);
  or OR_14812(g11737,g8359,g8292);
  or OR_14813(g12768,g7785,g7202);
  or OR_14814(g12832,g10347,g10348);
  or OR_14815(g12911,g10278,g12768);
  or OR_14816(g12925,g8928,g10511);
  or OR_14817(g12954,g12186,g9906);
  or OR_14818(g12981,g12219,g9967);
  or OR_14819(g12982,g12220,g9968);
  or OR_14820(g13006,g12284,g10034);
  or OR_14821(g13077,g11330,g943);
  or OR_14822(g13091,g329,g319,g10796);
  or OR_14823(g13095,g11374,g1287);
  or OR_14824(g13155,g11496,g11546);
  or OR_14825(g13211,g11294,g7567);
  or OR_14826(g13242,g11336,g7601);
  or OR_14827(g13289,g10619,g10624);
  or OR_14828(g13295,g10625,g10655);
  or OR_14829(g13296,g10626,g10657);
  or OR_14830(g13300,g10656,g10676);
  or OR_14831(g13385,g11967,g9479);
  or OR_14832(g13526,g209,g10685,g301);
  or OR_14833(g13540,g10822,g10827);
  or OR_14834(g13543,g10543,g10565);
  or OR_14835(g13570,g9223,g11130);
  or OR_14836(g13597,g9247,g11149);
  or OR_14837(g13623,g482,g12527);
  or OR_14838(g13657,g7251,g10616);
  or OR_14839(g13660,g8183,g12527);
  or OR_14840(g13662,g10896,g10917);
  or OR_14841(g13699,g10921,g10947);
  or OR_14842(g13728,g6804,g12527);
  or OR_14843(g13761,g490,g12527);
  or OR_14844(g13762,g499,g12527);
  or OR_14845(g13794,g7396,g10684);
  or OR_14846(g13820,g11184,g9187,g12527);
  or OR_14847(g13858,g209,g10685);
  or OR_14848(g13888,g2941,g11691);
  or OR_14849(g13914,g8643,g11380);
  or OR_14850(g13938,g11213,g11191);
  or OR_14851(g13941,g11019,g11023);
  or OR_14852(g13969,g11448,g8913);
  or OR_14853(g13972,g11232,g11203);
  or OR_14854(g13973,g11024,g11028);
  or OR_14855(g13997,g11029,g11036);
  or OR_14856(g14030,g11037,g11046);
  or OR_14857(g14044,g10776,g8703);
  or OR_14858(g14062,g11047,g11116);
  or OR_14859(g14078,g10776,g8703);
  or OR_14860(g14119,g10776,g8703);
  or OR_14861(g14182,g11741,g11721,g753);
  or OR_14862(g14187,g8871,g11771);
  or OR_14863(g14309,g10320,g11048);
  or OR_14864(g14387,g9086,g11048);
  or OR_14865(g14511,g10685,g546);
  or OR_14866(g14583,g10685,g542);
  or OR_14867(g14844,g10776,g8703);
  or OR_14868(g14888,g10776,g8703);
  or OR_14869(g14936,g10776,g8703);
  or OR_14870(g14977,g10776,g8703);
  or OR_14871(g15017,g10776,g8703);
  or OR_14872(g15124,g13605,g4581);
  or OR_14873(g15125,g10363,g13605);
  or OR_14874(g15582,g8977,g12925);
  or OR_14875(g15727,g13383,g13345,g13333,g11010);
  or OR_14876(g15732,g13411,g13384,g13349,g11016);
  or OR_14877(g15789,g10819,g13211);
  or OR_14878(g15792,g12920,g10501);
  or OR_14879(g15800,g10821,g13242);
  or OR_14880(g15803,g12924,g10528);
  or OR_14881(g15910,g13025,g10654);
  or OR_14882(g15935,g13029,g10665);
  or OR_14883(g15965,g13035,g10675);
  or OR_14884(g15968,g13038,g10677);
  or OR_14885(g16021,g13047,g10706);
  or OR_14886(g16022,g13048,g10707);
  or OR_14887(g16052,g13060,g10724);
  or OR_14888(g16076,g13081,g10736);
  or OR_14889(g16173,g8796,g13464);
  or OR_14890(g16187,g8822,g13486);
  or OR_14891(g16239,g7892,g13432);
  or OR_14892(g16258,g13247,g10856);
  or OR_14893(g16261,g7898,g13469);
  or OR_14894(g16430,g182,g13657);
  or OR_14895(g16448,g13287,g10934);
  or OR_14896(g16506,g13294,g10966);
  or OR_14897(g16800,g13436,g11027);
  or OR_14898(g16810,g13461,g11032);
  or OR_14899(g16811,g8690,g13914);
  or OR_14900(g16839,g13473,g11035);
  or OR_14901(g16866,g13492,g11044);
  or OR_14902(g16867,g13493,g11045);
  or OR_14903(g16876,g14028,g11773,g11755);
  or OR_14904(g16882,g13508,g11114);
  or OR_14905(g16883,g13509,g11115);
  or OR_14906(g16926,g14061,g11804,g11780);
  or OR_14907(g16927,g13524,g11126);
  or OR_14908(g16928,g13525,g11127);
  or OR_14909(g16959,g13542,g11142);
  or OR_14910(g16970,g13567,g11163);
  or OR_14911(g17264,g7118,g14309);
  or OR_14912(g17268,g9220,g14387);
  or OR_14913(I18385,g14413,g14391,g14360);
  or OR_14914(g17464,g14334,g14313,g11935,I18385);
  or OR_14915(I18417,g14444,g14414,g14392);
  or OR_14916(g17488,g14361,g14335,g11954,I18417);
  or OR_14917(I18421,g14447,g14417,g14395);
  or OR_14918(g17490,g14364,g14337,g11958,I18421);
  or OR_14919(I18449,g14512,g14445,g14415);
  or OR_14920(g17510,g14393,g14362,g11972,I18449);
  or OR_14921(I18452,g14514,g14448,g14418);
  or OR_14922(g17511,g14396,g14365,g11976,I18452);
  or OR_14923(I18492,g14538,g14513,g14446);
  or OR_14924(g17569,g14416,g14394,g11995,I18492);
  or OR_14925(I18495,g14539,g14515,g14449);
  or OR_14926(g17570,g14419,g14397,g11999,I18495);
  or OR_14927(I18543,g14568,g14540,g14516);
  or OR_14928(g17594,g14450,g14420,g12025,I18543);
  or OR_14929(g18879,g17365,g14423);
  or OR_14930(g18994,g16303,g13632);
  or OR_14931(g19267,g17752,g17768);
  or OR_14932(g19274,g17753,g14791);
  or OR_14933(g19336,g17769,g14831);
  or OR_14934(g19337,g17770,g17785);
  or OR_14935(g19344,g17771,g14832);
  or OR_14936(g19356,g17784,g14874);
  or OR_14937(g19359,g17786,g14875);
  or OR_14938(g19363,g17810,g14913);
  or OR_14939(g19441,g15507,g12931);
  or OR_14940(g19449,g15567,g12939);
  or OR_14941(g19467,g16896,g14097);
  or OR_14942(g19475,g16930,g14126);
  or OR_14943(g19486,g15589,g12979);
  or OR_14944(g19488,g16965,g14148);
  or OR_14945(g19501,g16986,g14168);
  or OR_14946(g19522,g17057,g14180);
  or OR_14947(g19525,g7696,g16811);
  or OR_14948(g19534,g15650,g13019);
  or OR_14949(g19535,g15651,g13020);
  or OR_14950(g19555,g15672,g13030);
  or OR_14951(g19557,g17123,g14190);
  or OR_14952(g19572,g17133,g14193);
  or OR_14953(g19575,g15693,g13042);
  or OR_14954(g19576,g17138,g14202);
  or OR_14955(g19587,g15700,g13046);
  or OR_14956(g19593,g17145,g14210);
  or OR_14957(g19595,g17149,g14218);
  or OR_14958(g19604,g15704,g13059);
  or OR_14959(g19605,g15707,g13063);
  or OR_14960(g19619,g15712,g13080);
  or OR_14961(g19879,g15841,g13265);
  or OR_14962(g19904,g17636,g14654);
  or OR_14963(g19949,g17671,g14681);
  or OR_14964(g20034,g15902,g13299);
  or OR_14965(g20051,g15936,g13306);
  or OR_14966(g20063,g15978,g13313);
  or OR_14967(g20077,g16025,g13320);
  or OR_14968(g20082,g16026,g13321);
  or OR_14969(g20083,g2902,g17058);
  or OR_14970(g20148,g16128,g13393);
  or OR_14971(g20160,g16163,g13415);
  or OR_14972(g20169,g16184,g13460);
  or OR_14973(g20187,g16202,g13491);
  or OR_14974(g20196,g16207,g13497);
  or OR_14975(g20202,g16211,g13507);
  or OR_14976(g20217,g16221,g13523);
  or OR_14977(g20241,g16233,g13541);
  or OR_14978(g20276,g16243,g13566);
  or OR_14979(g20522,g691,g16893);
  or OR_14980(g20905,g7216,g17264);
  or OR_14981(g21891,g19948,g15103);
  or OR_14982(g21892,g19788,g15104);
  or OR_14983(g21893,g20094,g18655);
  or OR_14984(g21894,g20112,g15107);
  or OR_14985(g21895,g20135,g15108);
  or OR_14986(g21896,g20084,g15110);
  or OR_14987(g21897,g20095,g15111);
  or OR_14988(g21898,g20152,g15112);
  or OR_14989(g21899,g20162,g15113);
  or OR_14990(g21900,g20977,g15114);
  or OR_14991(g21901,g21251,g15115);
  or OR_14992(g22152,g21188,g17469);
  or OR_14993(g22217,g21302,g17617);
  or OR_14994(g22225,g21332,g17654);
  or OR_14995(g22226,g21333,g17655);
  or OR_14996(g22304,g21347,g17693);
  or OR_14997(g22318,g21394,g17783);
  or OR_14998(g22331,g21405,g17809);
  or OR_14999(g22447,g21464,g12761);
  or OR_15000(g22487,g21512,g12794);
  or OR_15001(g22490,g21513,g12795);
  or OR_15002(g22516,g21559,g12817);
  or OR_15003(g22530,g16751,g20171);
  or OR_15004(g22531,g20773,g20922);
  or OR_15005(g22547,g16855,g20215);
  or OR_15006(g22585,g20915,g21061);
  or OR_15007(g22591,g18893,g18909);
  or OR_15008(g22625,g18910,g18933);
  or OR_15009(g22634,g18934,g15590);
  or OR_15010(g22636,g18943,g15611);
  or OR_15011(g22639,g18950,g15612);
  or OR_15012(g22640,g18951,g15613);
  or OR_15013(g22641,g18974,g15631);
  or OR_15014(g22644,g18981,g15632);
  or OR_15015(g22645,g18982,g15633);
  or OR_15016(g22648,g18987,g15652);
  or OR_15017(g22652,g18992,g15653);
  or OR_15018(g22653,g18993,g15654);
  or OR_15019(g22659,g19062,g15673);
  or OR_15020(g22662,g19069,g15679);
  or OR_15021(g22664,g19139,g15694);
  or OR_15022(g22669,g7763,g19525);
  or OR_15023(g22679,g19145,g15701);
  or OR_15024(g22684,g19206,g15703);
  or OR_15025(g22707,g20559,g17156);
  or OR_15026(g22708,g19266,g15711);
  or OR_15027(g22751,g19333,g15716);
  or OR_15028(g22832,g19354,g15722);
  or OR_15029(g22872,g19372,g19383);
  or OR_15030(g22901,g19384,g15745);
  or OR_15031(g23087,g19487,g15852);
  or OR_15032(g23129,g19500,g15863);
  or OR_15033(g23153,g19521,g15876);
  or OR_15034(I22267,g20236,g20133,g20111);
  or OR_15035(g23162,g20184,g20170,I22267);
  or OR_15036(g23171,g19536,g15903);
  or OR_15037(g23183,g19545,g15911);
  or OR_15038(I22280,g20271,g20150,g20134);
  or OR_15039(g23184,g20198,g20185,I22280);
  or OR_15040(g23193,g19556,g15937);
  or OR_15041(g23194,g19564,g19578);
  or OR_15042(g23197,g19571,g15966);
  or OR_15043(I22298,g20371,g20161,g20151);
  or OR_15044(g23198,g20214,g20199,I22298);
  or OR_15045(g23209,g19585,g19601);
  or OR_15046(g23217,g19588,g16023);
  or OR_15047(g23251,g19637,g16098);
  or OR_15048(g23255,g19655,g16122);
  or OR_15049(g23261,g19660,g16125);
  or OR_15050(g23262,g19661,g16126);
  or OR_15051(g23275,g19680,g16160);
  or OR_15052(g23276,g19681,g16161);
  or OR_15053(g23296,g19691,g16177);
  or OR_15054(g23297,g19692,g16178);
  or OR_15055(g23298,g19693,g16179);
  or OR_15056(g23317,g19715,g16191);
  or OR_15057(g23318,g19716,g16192);
  or OR_15058(g23319,g19717,g16193);
  or OR_15059(g23345,g19735,g16203);
  or OR_15060(g23346,g19736,g16204);
  or OR_15061(g23358,g19746,g16212);
  or OR_15062(g23374,g19767,g13514);
  or OR_15063(g23383,g19756,g16222);
  or OR_15064(g23405,g19791,g16245);
  or OR_15065(g23574,g20093,g20108);
  or OR_15066(g23615,g20109,g20131);
  or OR_15067(I22830,g21429,g21338,g21307);
  or OR_15068(g23687,g21384,g21363,I22830);
  or OR_15069(g23716,g9194,g20905);
  or OR_15070(g23720,g20165,g16801);
  or OR_15071(I22852,g21459,g21350,g21339);
  or OR_15072(g23721,g21401,g21385,I22852);
  or OR_15073(g23750,g20174,g16840);
  or OR_15074(I22880,g21509,g21356,g21351);
  or OR_15075(g23751,g21415,g21402,I22880);
  or OR_15076(g23770,g20188,g16868);
  or OR_15077(I22912,g21555,g21364,g21357);
  or OR_15078(g23771,g21432,g21416,I22912);
  or OR_15079(g23795,g20203,g16884);
  or OR_15080(I22958,g21603,g21386,g21365);
  or OR_15081(g23796,g21462,g21433,I22958);
  or OR_15082(g23822,g20218,g16929);
  or OR_15083(g23825,g20705,g20781);
  or OR_15084(g23989,g20581,g17179);
  or OR_15085(g23997,g20602,g17191);
  or OR_15086(I23162,g19919,g19968,g20014,g20841);
  or OR_15087(I23163,g20982,g21127,g21193,g21256);
  or OR_15088(g24151,g18088,g21661);
  or OR_15089(g24200,g22831,g18103);
  or OR_15090(g24201,g22848,g18104);
  or OR_15091(g24202,g22899,g18106);
  or OR_15092(g24203,g22982,g18107);
  or OR_15093(g24204,g22990,g18108);
  or OR_15094(g24205,g23006,g18109);
  or OR_15095(g24206,g23386,g18110);
  or OR_15096(g24207,g23396,g18119);
  or OR_15097(g24208,g23404,g18121);
  or OR_15098(g24209,g23415,g18122);
  or OR_15099(g24210,g22900,g18125);
  or OR_15100(g24211,g23572,g18138);
  or OR_15101(g24212,g23280,g18155);
  or OR_15102(g24213,g23220,g18186);
  or OR_15103(g24214,g23471,g18195);
  or OR_15104(g24215,g23484,g18196);
  or OR_15105(g24216,g23416,g18197);
  or OR_15106(g24231,g22589,g18201);
  or OR_15107(g24232,g22686,g18228);
  or OR_15108(g24233,g22590,g18236);
  or OR_15109(g24234,g22622,g18237);
  or OR_15110(g24235,g22632,g18238);
  or OR_15111(g24236,g22489,g18241);
  or OR_15112(g24237,g22515,g18242);
  or OR_15113(g24238,g23254,g18248);
  or OR_15114(g24239,g22752,g18250);
  or OR_15115(g24240,g22861,g18251);
  or OR_15116(g24241,g22920,g18252);
  or OR_15117(g24242,g22834,g18253);
  or OR_15118(g24243,g22992,g18254);
  or OR_15119(g24244,g23349,g18255);
  or OR_15120(g24245,g22849,g18256);
  or OR_15121(g24246,g23372,g18257);
  or OR_15122(g24247,g22623,g18259);
  or OR_15123(g24248,g22710,g18286);
  or OR_15124(g24249,g22624,g18294);
  or OR_15125(g24250,g22633,g18295);
  or OR_15126(g24251,g22637,g18296);
  or OR_15127(g24252,g22518,g18299);
  or OR_15128(g24253,g22525,g18300);
  or OR_15129(g24254,g23265,g18306);
  or OR_15130(g24255,g22835,g18308);
  or OR_15131(g24256,g22873,g18309);
  or OR_15132(g24257,g22938,g18310);
  or OR_15133(g24258,g22851,g18311);
  or OR_15134(g24259,g23008,g18312);
  or OR_15135(g24260,g23373,g18313);
  or OR_15136(g24261,g22862,g18314);
  or OR_15137(g24262,g23387,g18315);
  or OR_15138(g24263,g23497,g18529);
  or OR_15139(g24264,g22310,g18559);
  or OR_15140(g24265,g22316,g18560);
  or OR_15141(g24266,g22329,g18561);
  or OR_15142(g24267,g23439,g18611);
  or OR_15143(g24268,g23025,g18612);
  or OR_15144(g24269,g23131,g18613);
  or OR_15145(g24270,g23165,g18614);
  or OR_15146(g24271,g23451,g18628);
  or OR_15147(g24272,g23056,g18629);
  or OR_15148(g24273,g23166,g18630);
  or OR_15149(g24274,g23187,g18631);
  or OR_15150(g24275,g23474,g18645);
  or OR_15151(g24276,g23083,g18646);
  or OR_15152(g24277,g23188,g18647);
  or OR_15153(g24278,g23201,g18648);
  or OR_15154(g24279,g23218,g15105);
  or OR_15155(g24280,g23292,g15109);
  or OR_15156(g24281,g23397,g18656);
  or OR_15157(g24282,g23407,g18657);
  or OR_15158(g24334,g23991,g18676);
  or OR_15159(g24335,g22165,g18678);
  or OR_15160(g24336,g24012,g18753);
  or OR_15161(g24337,g23540,g18754);
  or OR_15162(g24338,g23658,g18755);
  or OR_15163(g24339,g23690,g18756);
  or OR_15164(g24340,g24016,g18770);
  or OR_15165(g24341,g23564,g18771);
  or OR_15166(g24342,g23691,g18772);
  or OR_15167(g24343,g23724,g18773);
  or OR_15168(g24344,g22145,g18787);
  or OR_15169(g24345,g23606,g18788);
  or OR_15170(g24346,g23725,g18789);
  or OR_15171(g24347,g23754,g18790);
  or OR_15172(g24348,g22149,g18804);
  or OR_15173(g24349,g23646,g18805);
  or OR_15174(g24350,g23755,g18806);
  or OR_15175(g24351,g23774,g18807);
  or OR_15176(g24352,g22157,g18821);
  or OR_15177(g24353,g23682,g18822);
  or OR_15178(g24354,g23775,g18823);
  or OR_15179(g24355,g23799,g18824);
  or OR_15180(g24363,g7831,g22138);
  or OR_15181(g24374,g19345,g24004);
  or OR_15182(g24390,g23779,g21285);
  or OR_15183(g24398,g23801,g21296);
  or OR_15184(g24401,g23811,g21298);
  or OR_15185(g24430,g23151,g8234);
  or OR_15186(g24432,g23900,g21361);
  or OR_15187(g24433,g10878,g22400);
  or OR_15188(g24443,g23917,g21378);
  or OR_15189(g24444,g10890,g22400);
  or OR_15190(g24447,g10948,g22450);
  or OR_15191(g24457,g10902,g22400);
  or OR_15192(g24460,g10967,g22450);
  or OR_15193(g24468,g10925,g22400);
  or OR_15194(g24471,g10999,g22450);
  or OR_15195(g24478,g11003,g22450);
  or OR_15196(g24496,g24008,g21557);
  or OR_15197(g24500,g24011,g21605);
  or OR_15198(g24510,g22488,g7567);
  or OR_15199(g24517,g22158,g18906);
  or OR_15200(g24518,g22517,g7601);
  or OR_15201(g24557,g22308,g19207);
  or OR_15202(I23755,g22904,g22927,g22980,g23444);
  or OR_15203(I23756,g23457,g23480,g23494,g23511);
  or OR_15204(g24561,I23755,I23756);
  or OR_15205(g24565,g22309,g19275);
  or OR_15206(g24577,g2856,g22531);
  or OR_15207(g24578,g2882,g23825);
  or OR_15208(g24580,g22340,g13096);
  or OR_15209(g24641,g22151,g22159);
  or OR_15210(g24653,g2848,g22585);
  or OR_15211(g24705,g2890,g23267);
  or OR_15212(g24715,g22189,g22207);
  or OR_15213(g24746,g22588,g19461);
  or OR_15214(g24782,g23857,g23872);
  or OR_15215(g24799,g23901,g23921);
  or OR_15216(g24813,g22685,g19594);
  or OR_15217(g24821,g21404,g23990);
  or OR_15218(g24840,g21419,g23996);
  or OR_15219(g24841,g21420,g23998);
  or OR_15220(g24842,g7804,g22669);
  or OR_15221(g24853,g21452,g24001);
  or OR_15222(g24854,g21453,g24002);
  or OR_15223(g24879,g21465,g24009);
  or OR_15224(g24896,g22863,g19684);
  or OR_15225(g24907,g21558,g24015);
  or OR_15226(g24919,g21606,g22143);
  or OR_15227(g24935,g22937,g19749);
  or OR_15228(g24946,g22360,g22409,g8130);
  or OR_15229(I24117,g23088,g23154,g23172);
  or OR_15230(g24952,g21326,g21340,I24117);
  or OR_15231(g24965,g22667,g23825);
  or OR_15232(g24968,g22360,g22409,g23389);
  or OR_15233(g25010,g23267,g2932);
  or OR_15234(g25037,g23103,g19911);
  or OR_15235(g25261,g23348,g20193);
  or OR_15236(g25539,g23531,g20628);
  or OR_15237(g25545,g23551,g20658);
  or OR_15238(g25575,g24139,g24140);
  or OR_15239(g25576,g24141,g24142);
  or OR_15240(g25577,g24143,g24144);
  or OR_15241(g25582,g21662,g24152);
  or OR_15242(g25583,g21666,g24153);
  or OR_15243(g25584,g21670,g24154);
  or OR_15244(g25585,g21674,g24155);
  or OR_15245(g25586,g21678,g24156);
  or OR_15246(g25587,g21682,g24157);
  or OR_15247(g25588,g21686,g24158);
  or OR_15248(g25589,g21690,g24159);
  or OR_15249(g25590,g21694,g24160);
  or OR_15250(g25591,g24642,g21705);
  or OR_15251(g25592,g24672,g21706);
  or OR_15252(g25593,g24716,g21707);
  or OR_15253(g25594,g24772,g21708);
  or OR_15254(g25595,g24835,g21717);
  or OR_15255(g25596,g24865,g21718);
  or OR_15256(g25597,g24892,g21719);
  or OR_15257(g25598,g24904,g21720);
  or OR_15258(g25599,g24914,g21721);
  or OR_15259(g25600,g24650,g18111);
  or OR_15260(g25601,g24660,g18112);
  or OR_15261(g25602,g24673,g18113);
  or OR_15262(g25603,g24698,g18114);
  or OR_15263(g25604,g24717,g18115);
  or OR_15264(g25605,g24743,g18116);
  or OR_15265(g25606,g24761,g18117);
  or OR_15266(g25607,g24773,g18118);
  or OR_15267(g25608,g24643,g18120);
  or OR_15268(g25609,g24915,g18126);
  or OR_15269(g25610,g24923,g18127);
  or OR_15270(g25611,g24931,g18128);
  or OR_15271(g25612,g24941,g18132);
  or OR_15272(g25613,g25181,g18140);
  or OR_15273(g25614,g24797,g18161);
  or OR_15274(g25615,g24803,g18162);
  or OR_15275(g25616,g25096,g18172);
  or OR_15276(g25617,g25466,g18189);
  or OR_15277(g25618,g25491,g18192);
  or OR_15278(g25619,g24961,g18193);
  or OR_15279(g25621,g24523,g18205);
  or OR_15280(g25622,g24546,g18217);
  or OR_15281(g25623,g24552,g18219);
  or OR_15282(g25624,g24408,g18224);
  or OR_15283(g25625,g24553,g18226);
  or OR_15284(g25626,g24499,g18235);
  or OR_15285(g25627,g24503,g18247);
  or OR_15286(g25628,g24600,g18249);
  or OR_15287(g25629,g24962,g18258);
  or OR_15288(g25630,g24532,g18263);
  or OR_15289(g25631,g24554,g18275);
  or OR_15290(g25632,g24558,g18277);
  or OR_15291(g25633,g24420,g18282);
  or OR_15292(g25634,g24559,g18284);
  or OR_15293(g25635,g24504,g18293);
  or OR_15294(g25636,g24507,g18305);
  or OR_15295(g25637,g24618,g18307);
  or OR_15296(g25638,g24977,g18316);
  or OR_15297(g25639,g25122,g18530);
  or OR_15298(g25643,g24602,g21736);
  or OR_15299(g25644,g24622,g21737);
  or OR_15300(g25645,g24679,g21738);
  or OR_15301(g25646,g24706,g21739);
  or OR_15302(g25647,g24725,g21740);
  or OR_15303(g25648,g24644,g21741);
  or OR_15304(g25649,g24654,g21742);
  or OR_15305(g25650,g24663,g21743);
  or OR_15306(g25651,g24680,g21744);
  or OR_15307(g25652,g24777,g21747);
  or OR_15308(g25653,g24664,g18602);
  or OR_15309(g25654,g24634,g18606);
  or OR_15310(g25655,g24645,g18607);
  or OR_15311(g25656,g24945,g18609);
  or OR_15312(g25657,g24624,g21782);
  or OR_15313(g25658,g24635,g21783);
  or OR_15314(g25659,g24707,g21784);
  or OR_15315(g25660,g24726,g21785);
  or OR_15316(g25661,g24754,g21786);
  or OR_15317(g25662,g24656,g21787);
  or OR_15318(g25663,g24666,g21788);
  or OR_15319(g25664,g24681,g21789);
  or OR_15320(g25665,g24708,g21790);
  or OR_15321(g25666,g24788,g21793);
  or OR_15322(g25667,g24682,g18619);
  or OR_15323(g25668,g24646,g18623);
  or OR_15324(g25669,g24657,g18624);
  or OR_15325(g25670,g24967,g18626);
  or OR_15326(g25671,g24637,g21828);
  or OR_15327(g25672,g24647,g21829);
  or OR_15328(g25673,g24727,g21830);
  or OR_15329(g25674,g24755,g21831);
  or OR_15330(g25675,g24769,g21832);
  or OR_15331(g25676,g24668,g21833);
  or OR_15332(g25677,g24684,g21834);
  or OR_15333(g25678,g24709,g21835);
  or OR_15334(g25679,g24728,g21836);
  or OR_15335(g25680,g24794,g21839);
  or OR_15336(g25681,g24710,g18636);
  or OR_15337(g25682,g24658,g18640);
  or OR_15338(g25683,g24669,g18641);
  or OR_15339(g25684,g24983,g18643);
  or OR_15340(g25685,g24476,g21866);
  or OR_15341(g25686,g24712,g21881);
  or OR_15342(g25687,g24729,g21882);
  or OR_15343(g25688,g24812,g21887);
  or OR_15344(g25689,g24849,g21888);
  or OR_15345(g25690,g24864,g21889);
  or OR_15346(g25691,g24536,g21890);
  or OR_15347(g25693,g24627,g18707);
  or OR_15348(g25694,g24638,g18738);
  or OR_15349(g25695,g24998,g21914);
  or OR_15350(g25696,g25012,g21915);
  or OR_15351(g25697,g25086,g21916);
  or OR_15352(g25698,g25104,g21917);
  or OR_15353(g25699,g25125,g21918);
  or OR_15354(g25700,g25040,g21919);
  or OR_15355(g25701,g25054,g21920);
  or OR_15356(g25702,g25068,g21921);
  or OR_15357(g25703,g25087,g21922);
  or OR_15358(g25704,g25173,g21925);
  or OR_15359(g25705,g25069,g18744);
  or OR_15360(g25706,g25030,g18748);
  or OR_15361(g25707,g25041,g18749);
  or OR_15362(g25708,g25526,g18751);
  or OR_15363(g25709,g25014,g21960);
  or OR_15364(g25710,g25031,g21961);
  or OR_15365(g25711,g25105,g21962);
  or OR_15366(g25712,g25126,g21963);
  or OR_15367(g25713,g25147,g21964);
  or OR_15368(g25714,g25056,g21965);
  or OR_15369(g25715,g25071,g21966);
  or OR_15370(g25716,g25088,g21967);
  or OR_15371(g25717,g25106,g21968);
  or OR_15372(g25718,g25187,g21971);
  or OR_15373(g25719,g25089,g18761);
  or OR_15374(g25720,g25042,g18765);
  or OR_15375(g25721,g25057,g18766);
  or OR_15376(g25722,g25530,g18768);
  or OR_15377(g25723,g25033,g22006);
  or OR_15378(g25724,g25043,g22007);
  or OR_15379(g25725,g25127,g22008);
  or OR_15380(g25726,g25148,g22009);
  or OR_15381(g25727,g25163,g22010);
  or OR_15382(g25728,g25076,g22011);
  or OR_15383(g25729,g25091,g22012);
  or OR_15384(g25730,g25107,g22013);
  or OR_15385(g25731,g25128,g22014);
  or OR_15386(g25732,g25201,g22017);
  or OR_15387(g25733,g25108,g18778);
  or OR_15388(g25734,g25058,g18782);
  or OR_15389(g25735,g25077,g18783);
  or OR_15390(g25736,g25536,g18785);
  or OR_15391(g25737,g25045,g22052);
  or OR_15392(g25738,g25059,g22053);
  or OR_15393(g25739,g25149,g22054);
  or OR_15394(g25740,g25164,g22055);
  or OR_15395(g25741,g25178,g22056);
  or OR_15396(g25742,g25093,g22057);
  or OR_15397(g25743,g25110,g22058);
  or OR_15398(g25744,g25129,g22059);
  or OR_15399(g25745,g25150,g22060);
  or OR_15400(g25746,g25217,g22063);
  or OR_15401(g25747,g25130,g18795);
  or OR_15402(g25748,g25078,g18799);
  or OR_15403(g25749,g25094,g18800);
  or OR_15404(g25750,g25543,g18802);
  or OR_15405(g25751,g25061,g22098);
  or OR_15406(g25752,g25079,g22099);
  or OR_15407(g25753,g25165,g22100);
  or OR_15408(g25754,g25179,g22101);
  or OR_15409(g25755,g25192,g22102);
  or OR_15410(g25756,g25112,g22103);
  or OR_15411(g25757,g25132,g22104);
  or OR_15412(g25758,g25151,g22105);
  or OR_15413(g25759,g25166,g22106);
  or OR_15414(g25760,g25238,g22109);
  or OR_15415(g25761,g25152,g18812);
  or OR_15416(g25762,g25095,g18816);
  or OR_15417(g25763,g25113,g18817);
  or OR_15418(g25764,g25551,g18819);
  or OR_15419(g25767,g25207,g12015);
  or OR_15420(g25774,g25223,g12043);
  or OR_15421(g25789,g25285,g14543);
  or OR_15422(g25791,g25411,g25371,g25328,g25290);
  or OR_15423(g25805,g25453,g25414,g25374,g25331);
  or OR_15424(g25819,g25323,g23836);
  or OR_15425(g25821,g25482,g25456,g25417,g25377);
  or OR_15426(g25834,g25366,g23854);
  or OR_15427(g25835,g25367,g23855);
  or OR_15428(g25836,g25368,g23856);
  or OR_15429(g25839,g25507,g25485,g25459,g25420);
  or OR_15430(g25856,g25518,g25510,g25488,g25462);
  or OR_15431(g25867,g25449,g23884);
  or OR_15432(g25868,g25450,g23885);
  or OR_15433(g25877,g25502,g23919);
  or OR_15434(g25878,g25503,g23920);
  or OR_15435(g25885,g25522,g23957);
  or OR_15436(g25894,g24817,g23229);
  or OR_15437(g25906,g25559,g24014);
  or OR_15438(g25910,g25565,g22142);
  or OR_15439(g25911,g22514,g24510);
  or OR_15440(g25917,g22524,g24518);
  or OR_15441(g25929,g24395,g22193);
  or OR_15442(g25935,g24402,g22208);
  or OR_15443(g25936,g24403,g22209);
  or OR_15444(g25937,g24406,g22216);
  or OR_15445(g25940,g24415,g22218);
  or OR_15446(g25941,g24416,g22219);
  or OR_15447(g25942,g24422,g22298);
  or OR_15448(g25943,g24423,g22299);
  or OR_15449(g25945,g24427,g22307);
  or OR_15450(g25960,g24566,g24678);
  or OR_15451(g26080,g19393,g24502);
  or OR_15452(g26082,g2898,g24561);
  or OR_15453(g26089,g24501,g22534);
  or OR_15454(g26099,g24506,g22538);
  or OR_15455(g26278,g24545,g24549);
  or OR_15456(g26293,g24550,g24555);
  or OR_15457(g26299,g24551,g22665);
  or OR_15458(g26305,g24556,g24564);
  or OR_15459(g26327,g8462,g24591);
  or OR_15460(g26328,g1183,g24591);
  or OR_15461(g26329,g8526,g24609);
  or OR_15462(g26334,g1171,g24591);
  or OR_15463(g26335,g1526,g24609);
  or OR_15464(g26342,g8407,g24591);
  or OR_15465(g26343,g1514,g24609);
  or OR_15466(g26344,g2927,g25010);
  or OR_15467(g26348,g8466,g24609);
  or OR_15468(g26349,g24630,g13409);
  or OR_15469(g26359,g24651,g22939);
  or OR_15470(g26361,g24674,g22991);
  or OR_15471(g26363,g2965,g24965);
  or OR_15472(g26365,g25504,g25141);
  or OR_15473(g26377,g24700,g23007);
  or OR_15474(g26386,g24719,g23023);
  or OR_15475(g26392,g24745,g23050);
  or OR_15476(g26396,g24762,g23062);
  or OR_15477(g26422,g24774,g23104);
  or OR_15478(g26512,g24786,g23130);
  or OR_15479(g26616,g24881,g24855,g24843,g24822);
  or OR_15480(g26636,g24897,g24884,g24858,g24846);
  or OR_15481(g26657,g24908,g24900,g24887,g24861);
  or OR_15482(g26673,g24433,g10674);
  or OR_15483(g26690,g10776,g24433);
  or OR_15484(g26694,g24444,g10704);
  or OR_15485(g26703,g24447,g10705);
  or OR_15486(g26721,g10776,g24444);
  or OR_15487(g26725,g24457,g10719);
  or OR_15488(g26733,g10776,g24447);
  or OR_15489(g26737,g24460,g10720);
  or OR_15490(g26751,g24903,g24912);
  or OR_15491(g26755,g10776,g24457);
  or OR_15492(g26759,g24468,g7511);
  or OR_15493(g26766,g10776,g24460);
  or OR_15494(g26770,g24471,g10732);
  or OR_15495(g26781,g24913,g24921);
  or OR_15496(g26785,g10776,g24468);
  or OR_15497(g26789,g10776,g24471);
  or OR_15498(g26793,g24478,g7520);
  or OR_15499(g26800,g24922,g24929);
  or OR_15500(g26805,g10776,g24478);
  or OR_15501(g26809,g24930,g24939);
  or OR_15502(g26813,g24940,g24949);
  or OR_15503(g26866,g20204,g20242,g24363);
  or OR_15504(I25612,g25567,g25568,g25569,g25570);
  or OR_15505(I25613,g25571,g25572,g25573,g25574);
  or OR_15506(g26874,I25612,I25613);
  or OR_15507(g26875,g21652,g25575);
  or OR_15508(g26876,g21655,g25576);
  or OR_15509(g26877,g21658,g25577);
  or OR_15510(g26878,g25578,g25579);
  or OR_15511(g26879,g25580,g25581);
  or OR_15512(g26880,g26610,g24186);
  or OR_15513(g26881,g26629,g24187);
  or OR_15514(g26882,g26650,g24188);
  or OR_15515(g26883,g26670,g24189);
  or OR_15516(g26884,g26511,g24190);
  or OR_15517(g26885,g26541,g24191);
  or OR_15518(g26886,g26651,g24192);
  or OR_15519(g26887,g26542,g24193);
  or OR_15520(g26888,g26671,g24194);
  or OR_15521(g26889,g26689,g24195);
  or OR_15522(g26890,g26630,g24196);
  or OR_15523(g26891,g26652,g24197);
  or OR_15524(g26892,g26719,g24198);
  or OR_15525(g26893,g26753,g24199);
  or OR_15526(g26894,g25979,g18129);
  or OR_15527(g26895,g26783,g18148);
  or OR_15528(g26896,g26341,g18171);
  or OR_15529(g26897,g26611,g18176);
  or OR_15530(g26898,g26387,g18194);
  or OR_15531(g26899,g26844,g18199);
  or OR_15532(g26900,g26819,g24217);
  or OR_15533(g26901,g26362,g24218);
  or OR_15534(g26902,g26378,g24219);
  or OR_15535(g26903,g26388,g24220);
  or OR_15536(g26904,g26393,g24221);
  or OR_15537(g26905,g26397,g24222);
  or OR_15538(g26906,g26423,g24223);
  or OR_15539(g26907,g26513,g24224);
  or OR_15540(g26908,g26358,g24225);
  or OR_15541(g26909,g26543,g24227);
  or OR_15542(g26910,g26571,g24228);
  or OR_15543(g26911,g26612,g24230);
  or OR_15544(g26912,g25946,g18209);
  or OR_15545(g26913,g25848,g18225);
  or OR_15546(g26914,g25949,g18227);
  or OR_15547(g26915,g25900,g18230);
  or OR_15548(g26916,g25916,g18232);
  or OR_15549(g26917,g26122,g18233);
  or OR_15550(g26918,g25931,g18243);
  or OR_15551(g26919,g25951,g18267);
  or OR_15552(g26920,g25865,g18283);
  or OR_15553(g26921,g25955,g18285);
  or OR_15554(g26922,g25902,g18288);
  or OR_15555(g26923,g25923,g18290);
  or OR_15556(g26924,g26153,g18291);
  or OR_15557(g26925,g25939,g18301);
  or OR_15558(g26926,g26633,g18531);
  or OR_15559(g26927,g26711,g18539);
  or OR_15560(g26928,g26713,g18541);
  or OR_15561(g26929,g26635,g18543);
  or OR_15562(g26930,g26799,g18544);
  or OR_15563(g26931,g26778,g18547);
  or OR_15564(g26932,g26684,g18549);
  or OR_15565(g26933,g26808,g18551);
  or OR_15566(g26934,g26845,g18556);
  or OR_15567(g26938,g26186,g21883);
  or OR_15568(g26939,g25907,g21884);
  or OR_15569(g26940,g25908,g21886);
  or OR_15570(g26944,g26130,g18658);
  or OR_15571(g26945,g26379,g24283);
  or OR_15572(g26946,g26389,g24284);
  or OR_15573(g26947,g26394,g24285);
  or OR_15574(g26948,g26399,g24286);
  or OR_15575(g26949,g26356,g24287);
  or OR_15576(g26950,g26357,g24288);
  or OR_15577(g26951,g26390,g24289);
  or OR_15578(g26952,g26360,g24290);
  or OR_15579(g26953,g26486,g24291);
  or OR_15580(g26954,g26380,g24292);
  or OR_15581(g26955,g26391,g24293);
  or OR_15582(g26956,g26487,g24294);
  or OR_15583(g26957,g26517,g24295);
  or OR_15584(g26958,g26395,g24297);
  or OR_15585(g26959,g26381,g24299);
  or OR_15586(g26960,g26258,g24304);
  or OR_15587(g26961,g26280,g24306);
  or OR_15588(g26962,g26295,g24307);
  or OR_15589(g26963,g26306,g24308);
  or OR_15590(g26964,g26259,g24316);
  or OR_15591(g26965,g26336,g24317);
  or OR_15592(g26966,g26345,g24318);
  or OR_15593(g26967,g26350,g24319);
  or OR_15594(g26968,g26307,g24321);
  or OR_15595(g26969,g26313,g24329);
  or OR_15596(g26970,g26308,g24332);
  or OR_15597(g26971,g26325,g24333);
  or OR_15598(g26972,g26780,g25229);
  or OR_15599(I25736,g12,g22150,g20277);
  or OR_15600(g27008,g26866,g21370,I25736);
  or OR_15601(g27016,g26821,g14585);
  or OR_15602(g27019,g26822,g14610);
  or OR_15603(g27024,g26826,g17692);
  or OR_15604(g27026,g26828,g17726);
  or OR_15605(g27031,g26213,g26190,g26166,g26148);
  or OR_15606(g27037,g26236,g26218,g26195,g26171);
  or OR_15607(g27108,g22522,g25911);
  or OR_15608(g27122,g22537,g25917);
  or OR_15609(g27126,g24378,g25787);
  or OR_15610(g27133,g25788,g24392);
  or OR_15611(g27135,g24387,g25803);
  or OR_15612(g27147,g25802,g24399);
  or OR_15613(g27150,g25804,g24400);
  or OR_15614(g27152,g24393,g25817);
  or OR_15615(g27159,g25814,g12953);
  or OR_15616(g27179,g25816,g24409);
  or OR_15617(g27182,g25818,g24410);
  or OR_15618(g27205,g25833,g24421);
  or OR_15619(g27224,g25870,g15678);
  or OR_15620(g27225,g2975,g26364);
  or OR_15621(g27226,g25872,g24436);
  or OR_15622(g27231,g25873,g15699);
  or OR_15623(g27232,g25874,g24450);
  or OR_15624(g27233,g25876,g24451);
  or OR_15625(g27236,g24620,g25974);
  or OR_15626(g27238,g25879,g24464);
  or OR_15627(g27239,g25881,g24465);
  or OR_15628(g27240,g25883,g24467);
  or OR_15629(g27241,g24584,g25984);
  or OR_15630(g27243,g25884,g24475);
  or OR_15631(g27244,g24652,g25995);
  or OR_15632(g27248,g24880,g25953);
  or OR_15633(g27250,g25901,g15738);
  or OR_15634(g27253,g24661,g26052);
  or OR_15635(g27257,g25904,g24498);
  or OR_15636(g27258,g25905,g15749);
  or OR_15637(g27261,g24544,g25996);
  or OR_15638(g27271,g24547,g26053);
  or OR_15639(g27274,g15779,g25915);
  or OR_15640(g27278,g15786,g25921);
  or OR_15641(g27283,g25922,g25924);
  or OR_15642(g27289,g25925,g25927);
  or OR_15643(g27290,g25926,g25928);
  or OR_15644(g27383,g24569,g25961);
  or OR_15645(g27394,g25957,g24573);
  or OR_15646(g27403,g25962,g24581);
  or OR_15647(g27405,g24572,g25968);
  or OR_15648(g27426,g25967,g24588);
  or OR_15649(g27429,g25969,g24589);
  or OR_15650(g27431,g24582,g25977);
  or OR_15651(g27450,g2917,g26483);
  or OR_15652(g27453,g25976,g24606);
  or OR_15653(g27456,g25978,g24607);
  or OR_15654(g27458,g24590,g25989);
  or OR_15655(g27484,g25988,g24628);
  or OR_15656(g27487,g25990,g24629);
  or OR_15657(g27489,g24608,g26022);
  or OR_15658(g27506,g26021,g24639);
  or OR_15659(g27509,g26023,g24640);
  or OR_15660(g27515,g26051,g13431);
  or OR_15661(g27524,g26050,g24649);
  or OR_15662(g27532,g16176,g26084);
  or OR_15663(g27533,g26078,g24659);
  or OR_15664(g27542,g16190,g26094);
  or OR_15665(g27543,g26085,g24670);
  or OR_15666(g27544,g26087,g24671);
  or OR_15667(g27551,g26091,g24675);
  or OR_15668(g27552,g26092,g24676);
  or OR_15669(g27555,g26095,g24686);
  or OR_15670(g27556,g26097,g24687);
  or OR_15671(g27561,g26100,g24702);
  or OR_15672(g27562,g26102,g24703);
  or OR_15673(g27563,g26104,g24704);
  or OR_15674(g27566,g26119,g24713);
  or OR_15675(g27567,g26121,g24714);
  or OR_15676(g27569,g26124,g24721);
  or OR_15677(g27570,g26126,g24722);
  or OR_15678(g27571,g26127,g24723);
  or OR_15679(g27572,g26129,g24724);
  or OR_15680(g27574,g26145,g24730);
  or OR_15681(g27575,g26147,g24731);
  or OR_15682(g27578,g26155,g24747);
  or OR_15683(g27579,g26157,g24748);
  or OR_15684(g27580,g26159,g24749);
  or OR_15685(g27581,g26161,g24750);
  or OR_15686(g27584,g26165,g24758);
  or OR_15687(g27589,g26177,g24763);
  or OR_15688(g27590,g26179,g24764);
  or OR_15689(g27591,g26181,g24765);
  or OR_15690(g27596,g26207,g24775);
  or OR_15691(g27663,g26323,g24820);
  or OR_15692(g27742,g17292,g26673);
  or OR_15693(g27779,g17317,g26694);
  or OR_15694(g27800,g17321,g26703);
  or OR_15695(g27837,g17401,g26725);
  or OR_15696(g27858,g17405,g26737);
  or OR_15697(g27886,g14438,g26759);
  or OR_15698(g27907,g17424,g26770);
  or OR_15699(g27937,g14506,g26793);
  or OR_15700(g27970,g26514,g25050);
  or OR_15701(g27972,g26131,g26105);
  or OR_15702(g27974,g26544,g25063);
  or OR_15703(g27980,g26105,g26131);
  or OR_15704(g28030,g24018,g26874);
  or OR_15705(I26522,g19890,g19935,g19984,g26365);
  or OR_15706(I26523,g20720,g20857,g20998,g21143);
  or OR_15707(g28041,g24145,g26878);
  or OR_15708(g28042,g24148,g26879);
  or OR_15709(g28043,g27323,g21714);
  or OR_15710(g28044,g27256,g18130);
  or OR_15711(g28045,g27378,g18141);
  or OR_15712(g28046,g27667,g18157);
  or OR_15713(g28047,g27676,g18160);
  or OR_15714(g28048,g27362,g18163);
  or OR_15715(g28049,g27684,g18164);
  or OR_15716(g28050,g27692,g18165);
  or OR_15717(g28051,g27699,g18166);
  or OR_15718(g28052,g27710,g18167);
  or OR_15719(g28053,g27393,g18168);
  or OR_15720(g28054,g27723,g18170);
  or OR_15721(g28055,g27560,g18190);
  or OR_15722(g28056,g27230,g18210);
  or OR_15723(g28057,g27033,g18218);
  or OR_15724(g28058,g27235,g18268);
  or OR_15725(g28059,g27042,g18276);
  or OR_15726(g28060,g27616,g18532);
  or OR_15727(g28061,g27287,g21735);
  or OR_15728(g28062,g27288,g21746);
  or OR_15729(g28063,g27541,g21773);
  or OR_15730(g28064,g27298,g21781);
  or OR_15731(g28065,g27299,g21792);
  or OR_15732(g28066,g27553,g21819);
  or OR_15733(g28067,g27309,g21827);
  or OR_15734(g28068,g27310,g21838);
  or OR_15735(g28069,g27564,g21865);
  or OR_15736(g28070,g27050,g21867);
  or OR_15737(g28071,g27085,g21873);
  or OR_15738(g28072,g27086,g21874);
  or OR_15739(g28073,g27097,g21875);
  or OR_15740(g28074,g27119,g21876);
  or OR_15741(g28075,g27083,g21877);
  or OR_15742(g28076,g27098,g21878);
  or OR_15743(g28077,g27120,g21879);
  or OR_15744(g28078,g27140,g21880);
  or OR_15745(g28082,g27369,g24315);
  or OR_15746(g28083,g27249,g18689);
  or OR_15747(g28084,g27254,g18698);
  or OR_15748(g28085,g27263,g18700);
  or OR_15749(g28086,g27268,g18702);
  or OR_15750(g28087,g27255,g18720);
  or OR_15751(g28088,g27264,g18729);
  or OR_15752(g28089,g27269,g18731);
  or OR_15753(g28090,g27275,g18733);
  or OR_15754(g28091,g27665,g21913);
  or OR_15755(g28092,g27666,g21924);
  or OR_15756(g28093,g27981,g21951);
  or OR_15757(g28094,g27673,g21959);
  or OR_15758(g28095,g27674,g21970);
  or OR_15759(g28096,g27988,g21997);
  or OR_15760(g28097,g27682,g22005);
  or OR_15761(g28098,g27683,g22016);
  or OR_15762(g28099,g27992,g22043);
  or OR_15763(g28100,g27690,g22051);
  or OR_15764(g28101,g27691,g22062);
  or OR_15765(g28102,g27995,g22089);
  or OR_15766(g28103,g27696,g22097);
  or OR_15767(g28104,g27697,g22108);
  or OR_15768(g28105,g27997,g22135);
  or OR_15769(g28118,g27821,g26815);
  or OR_15770(g28132,g27932,g27957);
  or OR_15771(g28134,g27958,g27962);
  or OR_15772(g28135,g27959,g27963);
  or OR_15773(g28138,g27964,g27968);
  or OR_15774(I26643,g27073,g27058,g27045,g27040);
  or OR_15775(I26644,g27057,g27044,g27039,g27032);
  or OR_15776(g28140,I26643,I26644);
  or OR_15777(g28172,g27469,g27440,g27416,g27395);
  or OR_15778(g28179,g27494,g27474,g27445,g27421);
  or OR_15779(g28180,g20242,g27511);
  or OR_15780(g28186,g27209,g27185,g27161,g27146);
  or OR_15781(g28188,g22535,g27108);
  or OR_15782(g28191,g27217,g27210,g27186,g27162);
  or OR_15783(g28194,g22540,g27122);
  or OR_15784(g28208,g27025,g27028);
  or OR_15785(g28209,g27223,g27141);
  or OR_15786(g28211,g27029,g27034);
  or OR_15787(g28212,g27030,g27035);
  or OR_15788(g28216,g27036,g27043);
  or OR_15789(I26741,g22881,g22905,g22928,g27402);
  or OR_15790(I26742,g23430,g23445,g23458,g23481);
  or OR_15791(g28220,g23495,I26741,I26742);
  or OR_15792(g28230,g27669,g14261);
  or OR_15793(g28279,g27087,g25909);
  or OR_15794(g28286,g27090,g15757);
  or OR_15795(g28295,g27094,g15783);
  or OR_15796(g28296,g27095,g15784);
  or OR_15797(g28297,g27096,g15785);
  or OR_15798(g28305,g27103,g15793);
  or OR_15799(g28306,g27104,g15794);
  or OR_15800(g28308,g27105,g15795);
  or OR_15801(g28309,g27106,g15796);
  or OR_15802(g28310,g27107,g15797);
  or OR_15803(g28316,g27113,g15804);
  or OR_15804(g28317,g27114,g15805);
  or OR_15805(g28319,g27115,g15807);
  or OR_15806(g28320,g27116,g15808);
  or OR_15807(g28322,g27117,g15809);
  or OR_15808(g28323,g27118,g15810);
  or OR_15809(g28328,g27127,g15812);
  or OR_15810(g28329,g27128,g15813);
  or OR_15811(g28331,g27129,g15814);
  or OR_15812(g28332,g27130,g15815);
  or OR_15813(g28334,g27131,g15817);
  or OR_15814(g28335,g27132,g15818);
  or OR_15815(g28342,g27134,g15819);
  or OR_15816(g28344,g27136,g15820);
  or OR_15817(g28345,g27137,g15821);
  or OR_15818(g28347,g27138,g15822);
  or OR_15819(g28348,g27139,g15823);
  or OR_15820(g28357,g27148,g15836);
  or OR_15821(g28358,g27149,g15837);
  or OR_15822(g28359,g27151,g15838);
  or OR_15823(g28361,g27153,g15839);
  or OR_15824(g28362,g27154,g15840);
  or OR_15825(g28368,g27158,g27184);
  or OR_15826(g28369,g27160,g25938);
  or OR_15827(g28371,g27177,g15847);
  or OR_15828(g28372,g27178,g15848);
  or OR_15829(g28373,g27180,g15849);
  or OR_15830(g28374,g27181,g15850);
  or OR_15831(g28375,g27183,g15851);
  or OR_15832(g28385,g27201,g15857);
  or OR_15833(g28386,g27202,g13277);
  or OR_15834(g28387,g27203,g15858);
  or OR_15835(g28388,g27204,g15859);
  or OR_15836(g28389,g27206,g15860);
  or OR_15837(g28390,g27207,g15861);
  or OR_15838(g28400,g27211,g15870);
  or OR_15839(g28401,g27212,g15871);
  or OR_15840(g28402,g27213,g15873);
  or OR_15841(g28403,g27214,g13282);
  or OR_15842(g28404,g27215,g15874);
  or OR_15843(g28405,g27216,g15875);
  or OR_15844(g28416,g27218,g15880);
  or OR_15845(g28417,g27219,g15881);
  or OR_15846(g28418,g27220,g15882);
  or OR_15847(g28419,g27221,g15884);
  or OR_15848(g28420,g27222,g13290);
  or OR_15849(g28428,g27227,g15912);
  or OR_15850(g28429,g27228,g15913);
  or OR_15851(g28430,g27229,g15914);
  or OR_15852(g28435,g27234,g15967);
  or OR_15853(g28490,g27262,g16185);
  or OR_15854(g28497,g27267,g16199);
  or OR_15855(g28511,g27272,g16208);
  or OR_15856(g28513,g27276,g26123);
  or OR_15857(g28517,g27280,g26154);
  or OR_15858(g28518,g27281,g26158);
  or OR_15859(g28525,g27284,g26176);
  or OR_15860(g28526,g27285,g26178);
  or OR_15861(g28527,g27286,g26182);
  or OR_15862(g28533,g27291,g26203);
  or OR_15863(g28534,g27292,g26204);
  or OR_15864(g28536,g27293,g26205);
  or OR_15865(g28538,g27294,g26206);
  or OR_15866(g28544,g27300,g26229);
  or OR_15867(g28545,g27301,g26230);
  or OR_15868(g28546,g27302,g26231);
  or OR_15869(g28548,g27303,g26232);
  or OR_15870(g28549,g27304,g26233);
  or OR_15871(g28551,g27305,g26234);
  or OR_15872(g28560,g27311,g26249);
  or OR_15873(g28561,g27312,g26250);
  or OR_15874(g28562,g27313,g26251);
  or OR_15875(g28564,g27314,g26252);
  or OR_15876(g28565,g27315,g26253);
  or OR_15877(g28566,g27316,g26254);
  or OR_15878(g28574,g27324,g26270);
  or OR_15879(g28576,g27325,g26271);
  or OR_15880(g28577,g27326,g26272);
  or OR_15881(g28578,g27327,g26273);
  or OR_15882(g28580,g27328,g26275);
  or OR_15883(g28581,g27329,g26276);
  or OR_15884(g28582,g27330,g26277);
  or OR_15885(g28589,g27331,g26285);
  or OR_15886(g28591,g27332,g26286);
  or OR_15887(g28592,g27333,g26288);
  or OR_15888(g28594,g27334,g26289);
  or OR_15889(g28595,g27335,g26290);
  or OR_15890(g28596,g27336,g26291);
  or OR_15891(g28600,g27339,g16427);
  or OR_15892(g28603,g27340,g26300);
  or OR_15893(g28605,g27341,g26302);
  or OR_15894(g28607,g27342,g26303);
  or OR_15895(g28609,g27346,g16483);
  or OR_15896(g28610,g27347,g16484);
  or OR_15897(g28611,g27348,g16485);
  or OR_15898(g28613,g27350,g26310);
  or OR_15899(g28614,g27351,g26311);
  or OR_15900(g28618,g27357,g16516);
  or OR_15901(g28619,g27358,g16517);
  or OR_15902(g28621,g27359,g16518);
  or OR_15903(g28622,g27360,g16519);
  or OR_15904(g28623,g27361,g16520);
  or OR_15905(g28625,g27363,g26324);
  or OR_15906(g28628,g27370,g16531);
  or OR_15907(g28629,g27371,g16532);
  or OR_15908(g28631,g27372,g16534);
  or OR_15909(g28632,g27373,g16535);
  or OR_15910(g28634,g27374,g16536);
  or OR_15911(g28635,g27375,g16537);
  or OR_15912(g28636,g27376,g16538);
  or OR_15913(g28640,g27384,g16590);
  or OR_15914(g28641,g27385,g16591);
  or OR_15915(g28643,g27386,g16592);
  or OR_15916(g28644,g27387,g16593);
  or OR_15917(g28646,g27388,g16595);
  or OR_15918(g28647,g27389,g16596);
  or OR_15919(g28649,g27390,g16597);
  or OR_15920(g28650,g27391,g16598);
  or OR_15921(g28651,g27392,g16599);
  or OR_15922(g28659,g27404,g16610);
  or OR_15923(g28661,g27406,g16611);
  or OR_15924(g28662,g27407,g16612);
  or OR_15925(g28664,g27408,g16613);
  or OR_15926(g28665,g27409,g16614);
  or OR_15927(g28667,g27410,g16616);
  or OR_15928(g28668,g27411,g16617);
  or OR_15929(g28670,g27412,g16618);
  or OR_15930(g28671,g27413,g16619);
  or OR_15931(g28680,g27427,g16633);
  or OR_15932(g28681,g27428,g16634);
  or OR_15933(g28682,g27430,g16635);
  or OR_15934(g28684,g27432,g16636);
  or OR_15935(g28685,g27433,g16637);
  or OR_15936(g28687,g27434,g16638);
  or OR_15937(g28688,g27435,g16639);
  or OR_15938(g28690,g27436,g16641);
  or OR_15939(g28691,g27437,g16642);
  or OR_15940(g28698,g27451,g16666);
  or OR_15941(g28699,g27452,g16667);
  or OR_15942(g28700,g27454,g16668);
  or OR_15943(g28701,g27455,g16669);
  or OR_15944(g28702,g27457,g16670);
  or OR_15945(g28704,g27459,g16671);
  or OR_15946(g28705,g27460,g16672);
  or OR_15947(g28707,g27461,g16673);
  or OR_15948(g28708,g27462,g16674);
  or OR_15949(g28715,g27480,g16700);
  or OR_15950(g28716,g27481,g13887);
  or OR_15951(g28717,g27482,g16701);
  or OR_15952(g28718,g27483,g16702);
  or OR_15953(g28719,g27485,g16703);
  or OR_15954(g28720,g27486,g16704);
  or OR_15955(g28721,g27488,g16705);
  or OR_15956(g28723,g27490,g16706);
  or OR_15957(g28724,g27491,g16707);
  or OR_15958(g28727,g27500,g16729);
  or OR_15959(g28728,g27501,g16730);
  or OR_15960(g28729,g27502,g16732);
  or OR_15961(g28730,g27503,g13912);
  or OR_15962(g28731,g27504,g16733);
  or OR_15963(g28732,g27505,g16734);
  or OR_15964(g28733,g27507,g16735);
  or OR_15965(g28734,g27508,g16736);
  or OR_15966(g28735,g27510,g16737);
  or OR_15967(g28743,g27517,g16758);
  or OR_15968(g28744,g27518,g16759);
  or OR_15969(g28745,g27519,g16760);
  or OR_15970(g28746,g27520,g16762);
  or OR_15971(g28747,g27521,g13942);
  or OR_15972(g28748,g27522,g16763);
  or OR_15973(g28749,g27523,g16764);
  or OR_15974(g28750,g27525,g16765);
  or OR_15975(g28751,g27526,g16766);
  or OR_15976(g28772,g27534,g16802);
  or OR_15977(g28773,g27535,g16803);
  or OR_15978(g28774,g27536,g16804);
  or OR_15979(g28775,g27537,g16806);
  or OR_15980(g28776,g27538,g13974);
  or OR_15981(g28777,g27539,g16807);
  or OR_15982(g28778,g27540,g16808);
  or OR_15983(g28814,g27545,g16841);
  or OR_15984(g28815,g27546,g16842);
  or OR_15985(g28816,g27547,g16843);
  or OR_15986(g28817,g27548,g16845);
  or OR_15987(g28818,g27549,g13998);
  or OR_15988(g28850,g27557,g16869);
  or OR_15989(g28851,g27558,g16870);
  or OR_15990(g28852,g27559,g16871);
  or OR_15991(g28884,g27568,g16885);
  or OR_15992(g29068,g27628,g17119);
  or OR_15993(g29078,g27633,g26572);
  or OR_15994(g29105,g27645,g17134);
  or OR_15995(g29114,g27646,g26602);
  or OR_15996(g29143,g27650,g17146);
  or OR_15997(g29148,g27651,g26606);
  or OR_15998(g29166,g27653,g17153);
  or OR_15999(g29168,g27658,g26613);
  or OR_16000(g29176,g27661,g17177);
  or OR_16001(g29197,g27187,g27163);
  or OR_16002(g29222,g28252,g18105);
  or OR_16003(g29223,g28341,g18131);
  or OR_16004(g29224,g28919,g18156);
  or OR_16005(g29225,g28451,g18158);
  or OR_16006(g29226,g28455,g18159);
  or OR_16007(g29227,g28456,g18169);
  or OR_16008(g29228,g28426,g18173);
  or OR_16009(g29229,g28532,g18191);
  or OR_16010(g29230,g28107,g18202);
  or OR_16011(g29231,g28301,g18229);
  or OR_16012(g29232,g28183,g18231);
  or OR_16013(g29233,g28171,g18234);
  or OR_16014(g29234,g28415,g18239);
  or OR_16015(g29235,g28110,g18260);
  or OR_16016(g29236,g28313,g18287);
  or OR_16017(g29237,g28185,g18289);
  or OR_16018(g29238,g28178,g18292);
  or OR_16019(g29239,g28427,g18297);
  or OR_16020(g29240,g28655,g18328);
  or OR_16021(g29241,g28638,g18332);
  or OR_16022(g29242,g28674,g18354);
  or OR_16023(g29243,g28657,g18358);
  or OR_16024(g29244,g28692,g18380);
  or OR_16025(g29245,g28676,g18384);
  or OR_16026(g29246,g28710,g18406);
  or OR_16027(g29247,g28694,g18410);
  or OR_16028(g29248,g28677,g18434);
  or OR_16029(g29249,g28658,g18438);
  or OR_16030(g29250,g28695,g18460);
  or OR_16031(g29251,g28679,g18464);
  or OR_16032(g29252,g28712,g18486);
  or OR_16033(g29253,g28697,g18490);
  or OR_16034(g29254,g28725,g18512);
  or OR_16035(g29255,g28714,g18516);
  or OR_16036(g29256,g28597,g18533);
  or OR_16037(g29257,g28228,g18600);
  or OR_16038(g29258,g28238,g18601);
  or OR_16039(g29259,g28304,g18603);
  or OR_16040(g29260,g28315,g18604);
  or OR_16041(g29261,g28247,g18605);
  or OR_16042(g29262,g28327,g18608);
  or OR_16043(g29263,g28239,g18617);
  or OR_16044(g29264,g28248,g18618);
  or OR_16045(g29265,g28318,g18620);
  or OR_16046(g29266,g28330,g18621);
  or OR_16047(g29267,g28257,g18622);
  or OR_16048(g29268,g28343,g18625);
  or OR_16049(g29269,g28249,g18634);
  or OR_16050(g29270,g28258,g18635);
  or OR_16051(g29271,g28333,g18637);
  or OR_16052(g29272,g28346,g18638);
  or OR_16053(g29273,g28269,g18639);
  or OR_16054(g29274,g28360,g18642);
  or OR_16055(g29275,g28165,g21868);
  or OR_16056(g29276,g28616,g18709);
  or OR_16057(g29277,g28440,g18710);
  or OR_16058(g29278,g28626,g18740);
  or OR_16059(g29279,g28442,g18741);
  or OR_16060(g29280,g28530,g18742);
  or OR_16061(g29281,g28541,g18743);
  or OR_16062(g29282,g28617,g18745);
  or OR_16063(g29283,g28627,g18746);
  or OR_16064(g29284,g28554,g18747);
  or OR_16065(g29285,g28639,g18750);
  or OR_16066(g29286,g28542,g18759);
  or OR_16067(g29287,g28555,g18760);
  or OR_16068(g29288,g28630,g18762);
  or OR_16069(g29289,g28642,g18763);
  or OR_16070(g29290,g28569,g18764);
  or OR_16071(g29291,g28660,g18767);
  or OR_16072(g29292,g28556,g18776);
  or OR_16073(g29293,g28570,g18777);
  or OR_16074(g29294,g28645,g18779);
  or OR_16075(g29295,g28663,g18780);
  or OR_16076(g29296,g28586,g18781);
  or OR_16077(g29297,g28683,g18784);
  or OR_16078(g29298,g28571,g18793);
  or OR_16079(g29299,g28587,g18794);
  or OR_16080(g29300,g28666,g18796);
  or OR_16081(g29301,g28686,g18797);
  or OR_16082(g29302,g28601,g18798);
  or OR_16083(g29303,g28703,g18801);
  or OR_16084(g29304,g28588,g18810);
  or OR_16085(g29305,g28602,g18811);
  or OR_16086(g29306,g28689,g18813);
  or OR_16087(g29307,g28706,g18814);
  or OR_16088(g29308,g28612,g18815);
  or OR_16089(g29309,g28722,g18818);
  or OR_16090(g29313,g28284,g27270);
  or OR_16091(g29319,g28812,g14453);
  or OR_16092(g29325,g28813,g27820);
  or OR_16093(g29366,g13738,g28439);
  or OR_16094(g29373,g13832,g28453);
  or OR_16095(g29476,g28108,g28112);
  or OR_16096(g29478,g28111,g22160);
  or OR_16097(g29479,g28113,g28116);
  or OR_16098(g29480,g28115,g22172);
  or OR_16099(g29481,g28117,g28125);
  or OR_16100(g29482,g28524,g27588);
  or OR_16101(g29483,g25801,g28130);
  or OR_16102(g29484,g28124,g22191);
  or OR_16103(g29485,g28535,g27594);
  or OR_16104(g29486,g28537,g27595);
  or OR_16105(g29487,g25815,g28133);
  or OR_16106(g29488,g28547,g27600);
  or OR_16107(g29489,g28550,g27601);
  or OR_16108(g29490,g25832,g28136);
  or OR_16109(g29495,g28563,g27614);
  or OR_16110(g29496,g28567,g27615);
  or OR_16111(g29501,g28583,g27634);
  or OR_16112(g29502,g28139,g25871);
  or OR_16113(g29504,g28143,g25875);
  or OR_16114(g29506,g28148,g25880);
  or OR_16115(g29508,g28152,g27041);
  or OR_16116(g29520,g28291,g28281,g28264,g28254);
  or OR_16117(g29529,g28303,g28293,g28283,g28267);
  or OR_16118(g29539,g2864,g28220);
  or OR_16119(g29583,g28182,g27099);
  or OR_16120(g29643,g28192,g27145);
  or OR_16121(g29692,g28197,g10873);
  or OR_16122(g29706,g28198,g27208);
  or OR_16123(g29716,g28199,g15856);
  or OR_16124(g29717,g28200,g10883);
  or OR_16125(g29730,g28150,g28141);
  or OR_16126(g29734,g28201,g15872);
  or OR_16127(g29735,g28202,g10898);
  or OR_16128(g29741,g28205,g15883);
  or OR_16129(g29748,g28210,g28214);
  or OR_16130(g29753,g28213,g22720);
  or OR_16131(g29754,g28215,g28218);
  or OR_16132(g29756,g22717,g28223);
  or OR_16133(g29763,g28217,g22762);
  or OR_16134(g29764,g28219,g28226);
  or OR_16135(g29768,g22760,g28229);
  or OR_16136(g29775,g25966,g28232);
  or OR_16137(g29776,g28225,g22846);
  or OR_16138(g29777,g28227,g28234);
  or OR_16139(g29786,g22843,g28240);
  or OR_16140(g29790,g25975,g28242);
  or OR_16141(g29791,g28233,g22859);
  or OR_16142(g29792,g28235,g28244);
  or OR_16143(g29793,g28237,g27247);
  or OR_16144(g29801,g25987,g28251);
  or OR_16145(g29802,g28243,g22871);
  or OR_16146(g29813,g26020,g28261);
  or OR_16147(g29848,g28260,g26077);
  or OR_16148(g29849,g26049,g28273);
  or OR_16149(g29864,g28272,g26086);
  or OR_16150(g29879,g28289,g26096);
  or OR_16151(g29892,g28300,g26120);
  or OR_16152(g29904,g28312,g26146);
  or OR_16153(I28147,g2946,g24561,g28220);
  or OR_16154(g29914,g22531,g22585,I28147);
  or OR_16155(g30081,g28454,g11366);
  or OR_16156(g30092,g28466,g16699);
  or OR_16157(g30093,g28467,g11397);
  or OR_16158(g30103,g28477,g16731);
  or OR_16159(g30104,g28478,g11427);
  or OR_16160(g30114,g28488,g16761);
  or OR_16161(g30115,g28489,g11449);
  or OR_16162(g30127,g28494,g16805);
  or OR_16163(g30128,g28495,g11497);
  or OR_16164(g30141,g28499,g16844);
  or OR_16165(g30163,g23381,g28523);
  or OR_16166(g30176,g23392,g28531);
  or OR_16167(g30189,g23401,g28543);
  or OR_16168(g30201,g23412,g28557);
  or OR_16169(g30214,g23424,g28572);
  or OR_16170(g30270,g28624,g27664);
  or OR_16171(g30279,g28637,g27668);
  or OR_16172(g30286,g28191,g28186);
  or OR_16173(g30287,g28653,g27677);
  or OR_16174(g30291,g28672,g27685);
  or OR_16175(g30293,g28236,g27246);
  or OR_16176(g30298,g28245,g27251);
  or OR_16177(g30300,g28246,g27252);
  or OR_16178(g30304,g28255,g27259);
  or OR_16179(g30307,g28256,g27260);
  or OR_16180(g30311,g28265,g27265);
  or OR_16181(g30314,g28268,g27266);
  or OR_16182(I28566,g29201,g29202,g29203,g28035);
  or OR_16183(I28567,g29204,g29205,g29206,g29207);
  or OR_16184(g30317,g29208,I28566,I28567);
  or OR_16185(g30333,g29834,g21699);
  or OR_16186(g30334,g29837,g18143);
  or OR_16187(g30335,g29746,g18174);
  or OR_16188(g30336,g29324,g18203);
  or OR_16189(g30337,g29334,g18220);
  or OR_16190(g30338,g29613,g18240);
  or OR_16191(g30339,g29629,g18244);
  or OR_16192(g30340,g29377,g18245);
  or OR_16193(g30341,g29380,g18246);
  or OR_16194(g30342,g29330,g18261);
  or OR_16195(g30343,g29344,g18278);
  or OR_16196(g30344,g29630,g18298);
  or OR_16197(g30345,g29644,g18302);
  or OR_16198(g30346,g29381,g18303);
  or OR_16199(g30347,g29383,g18304);
  or OR_16200(g30348,g30083,g18329);
  or OR_16201(g30349,g30051,g18333);
  or OR_16202(g30350,g30118,g18334);
  or OR_16203(g30351,g30084,g18339);
  or OR_16204(g30352,g30094,g18340);
  or OR_16205(g30353,g30095,g18355);
  or OR_16206(g30354,g30064,g18359);
  or OR_16207(g30355,g30131,g18360);
  or OR_16208(g30356,g30096,g18365);
  or OR_16209(g30357,g30107,g18366);
  or OR_16210(g30358,g30108,g18381);
  or OR_16211(g30359,g30075,g18385);
  or OR_16212(g30360,g30145,g18386);
  or OR_16213(g30361,g30109,g18391);
  or OR_16214(g30362,g30120,g18392);
  or OR_16215(g30363,g30121,g18407);
  or OR_16216(g30364,g30086,g18411);
  or OR_16217(g30365,g30158,g18412);
  or OR_16218(g30366,g30122,g18417);
  or OR_16219(g30367,g30133,g18418);
  or OR_16220(g30368,g30098,g18435);
  or OR_16221(g30369,g30066,g18439);
  or OR_16222(g30370,g30135,g18440);
  or OR_16223(g30371,g30099,g18445);
  or OR_16224(g30372,g30110,g18446);
  or OR_16225(g30373,g30111,g18461);
  or OR_16226(g30374,g30078,g18465);
  or OR_16227(g30375,g30149,g18466);
  or OR_16228(g30376,g30112,g18471);
  or OR_16229(g30377,g30124,g18472);
  or OR_16230(g30378,g30125,g18487);
  or OR_16231(g30379,g30089,g18491);
  or OR_16232(g30380,g30161,g18492);
  or OR_16233(g30381,g30126,g18497);
  or OR_16234(g30382,g30137,g18498);
  or OR_16235(g30383,g30138,g18513);
  or OR_16236(g30384,g30101,g18517);
  or OR_16237(g30385,g30172,g18518);
  or OR_16238(g30386,g30139,g18523);
  or OR_16239(g30387,g30151,g18524);
  or OR_16240(g30388,g30023,g18534);
  or OR_16241(g30389,g29969,g18554);
  or OR_16242(g30390,g29985,g18555);
  or OR_16243(g30391,g30080,g18557);
  or OR_16244(g30392,g30091,g18558);
  or OR_16245(g30393,g29986,g21748);
  or OR_16246(g30394,g29805,g21753);
  or OR_16247(g30395,g29841,g21754);
  or OR_16248(g30396,g29856,g21755);
  or OR_16249(g30397,g29747,g21756);
  or OR_16250(g30398,g29749,g21757);
  or OR_16251(g30399,g29757,g21758);
  or OR_16252(g30400,g29766,g21759);
  or OR_16253(g30401,g29782,g21760);
  or OR_16254(g30402,g29871,g21761);
  or OR_16255(g30403,g29750,g21762);
  or OR_16256(g30404,g29758,g21763);
  or OR_16257(g30405,g29767,g21764);
  or OR_16258(g30406,g29783,g21765);
  or OR_16259(g30407,g29794,g21766);
  or OR_16260(g30408,g29806,g21767);
  or OR_16261(g30409,g29842,g21768);
  or OR_16262(g30410,g29857,g21769);
  or OR_16263(g30411,g29872,g21770);
  or OR_16264(g30412,g29885,g21771);
  or OR_16265(g30413,g30001,g21772);
  or OR_16266(g30414,g30002,g21794);
  or OR_16267(g30415,g29843,g21799);
  or OR_16268(g30416,g29858,g21800);
  or OR_16269(g30417,g29874,g21801);
  or OR_16270(g30418,g29751,g21802);
  or OR_16271(g30419,g29759,g21803);
  or OR_16272(g30420,g29769,g21804);
  or OR_16273(g30421,g29784,g21805);
  or OR_16274(g30422,g29795,g21806);
  or OR_16275(g30423,g29887,g21807);
  or OR_16276(g30424,g29760,g21808);
  or OR_16277(g30425,g29770,g21809);
  or OR_16278(g30426,g29785,g21810);
  or OR_16279(g30427,g29796,g21811);
  or OR_16280(g30428,g29807,g21812);
  or OR_16281(g30429,g29844,g21813);
  or OR_16282(g30430,g29859,g21814);
  or OR_16283(g30431,g29875,g21815);
  or OR_16284(g30432,g29888,g21816);
  or OR_16285(g30433,g29899,g21817);
  or OR_16286(g30434,g30024,g21818);
  or OR_16287(g30435,g30025,g21840);
  or OR_16288(g30436,g29860,g21845);
  or OR_16289(g30437,g29876,g21846);
  or OR_16290(g30438,g29890,g21847);
  or OR_16291(g30439,g29761,g21848);
  or OR_16292(g30440,g29771,g21849);
  or OR_16293(g30441,g29787,g21850);
  or OR_16294(g30442,g29797,g21851);
  or OR_16295(g30443,g29808,g21852);
  or OR_16296(g30444,g29901,g21853);
  or OR_16297(g30445,g29772,g21854);
  or OR_16298(g30446,g29788,g21855);
  or OR_16299(g30447,g29798,g21856);
  or OR_16300(g30448,g29809,g21857);
  or OR_16301(g30449,g29845,g21858);
  or OR_16302(g30450,g29861,g21859);
  or OR_16303(g30451,g29877,g21860);
  or OR_16304(g30452,g29891,g21861);
  or OR_16305(g30453,g29902,g21862);
  or OR_16306(g30454,g29909,g21863);
  or OR_16307(g30455,g30041,g21864);
  or OR_16308(g30456,g29378,g21869);
  or OR_16309(g30457,g29369,g21885);
  or OR_16310(g30458,g30005,g24330);
  or OR_16311(g30459,g29314,g21926);
  or OR_16312(g30460,g30207,g21931);
  or OR_16313(g30461,g30219,g21932);
  or OR_16314(g30462,g30228,g21933);
  or OR_16315(g30463,g30140,g21934);
  or OR_16316(g30464,g30152,g21935);
  or OR_16317(g30465,g30164,g21936);
  or OR_16318(g30466,g30174,g21937);
  or OR_16319(g30467,g30185,g21938);
  or OR_16320(g30468,g30238,g21939);
  or OR_16321(g30469,g30153,g21940);
  or OR_16322(g30470,g30165,g21941);
  or OR_16323(g30471,g30175,g21942);
  or OR_16324(g30472,g30186,g21943);
  or OR_16325(g30473,g30196,g21944);
  or OR_16326(g30474,g30208,g21945);
  or OR_16327(g30475,g30220,g21946);
  or OR_16328(g30476,g30229,g21947);
  or OR_16329(g30477,g30239,g21948);
  or OR_16330(g30478,g30248,g21949);
  or OR_16331(g30479,g29320,g21950);
  or OR_16332(g30480,g29321,g21972);
  or OR_16333(g30481,g30221,g21977);
  or OR_16334(g30482,g30230,g21978);
  or OR_16335(g30483,g30241,g21979);
  or OR_16336(g30484,g30154,g21980);
  or OR_16337(g30485,g30166,g21981);
  or OR_16338(g30486,g30177,g21982);
  or OR_16339(g30487,g30187,g21983);
  or OR_16340(g30488,g30197,g21984);
  or OR_16341(g30489,g30250,g21985);
  or OR_16342(g30490,g30167,g21986);
  or OR_16343(g30491,g30178,g21987);
  or OR_16344(g30492,g30188,g21988);
  or OR_16345(g30493,g30198,g21989);
  or OR_16346(g30494,g30209,g21990);
  or OR_16347(g30495,g30222,g21991);
  or OR_16348(g30496,g30231,g21992);
  or OR_16349(g30497,g30242,g21993);
  or OR_16350(g30498,g30251,g21994);
  or OR_16351(g30499,g30261,g21995);
  or OR_16352(g30500,g29326,g21996);
  or OR_16353(g30501,g29327,g22018);
  or OR_16354(g30502,g30232,g22023);
  or OR_16355(g30503,g30243,g22024);
  or OR_16356(g30504,g30253,g22025);
  or OR_16357(g30505,g30168,g22026);
  or OR_16358(g30506,g30179,g22027);
  or OR_16359(g30507,g30190,g22028);
  or OR_16360(g30508,g30199,g22029);
  or OR_16361(g30509,g30210,g22030);
  or OR_16362(g30510,g30263,g22031);
  or OR_16363(g30511,g30180,g22032);
  or OR_16364(g30512,g30191,g22033);
  or OR_16365(g30513,g30200,g22034);
  or OR_16366(g30514,g30211,g22035);
  or OR_16367(g30515,g30223,g22036);
  or OR_16368(g30516,g30233,g22037);
  or OR_16369(g30517,g30244,g22038);
  or OR_16370(g30518,g30254,g22039);
  or OR_16371(g30519,g30264,g22040);
  or OR_16372(g30520,g30272,g22041);
  or OR_16373(g30521,g29331,g22042);
  or OR_16374(g30522,g29332,g22064);
  or OR_16375(g30523,g30245,g22069);
  or OR_16376(g30524,g30255,g22070);
  or OR_16377(g30525,g30266,g22071);
  or OR_16378(g30526,g30181,g22072);
  or OR_16379(g30527,g30192,g22073);
  or OR_16380(g30528,g30202,g22074);
  or OR_16381(g30529,g30212,g22075);
  or OR_16382(g30530,g30224,g22076);
  or OR_16383(g30531,g30274,g22077);
  or OR_16384(g30532,g30193,g22078);
  or OR_16385(g30533,g30203,g22079);
  or OR_16386(g30534,g30213,g22080);
  or OR_16387(g30535,g30225,g22081);
  or OR_16388(g30536,g30234,g22082);
  or OR_16389(g30537,g30246,g22083);
  or OR_16390(g30538,g30256,g22084);
  or OR_16391(g30539,g30267,g22085);
  or OR_16392(g30540,g30275,g22086);
  or OR_16393(g30541,g30281,g22087);
  or OR_16394(g30542,g29337,g22088);
  or OR_16395(g30543,g29338,g22110);
  or OR_16396(g30544,g30257,g22115);
  or OR_16397(g30545,g30268,g22116);
  or OR_16398(g30546,g30277,g22117);
  or OR_16399(g30547,g30194,g22118);
  or OR_16400(g30548,g30204,g22119);
  or OR_16401(g30549,g30215,g22120);
  or OR_16402(g30550,g30226,g22121);
  or OR_16403(g30551,g30235,g22122);
  or OR_16404(g30552,g30283,g22123);
  or OR_16405(g30553,g30205,g22124);
  or OR_16406(g30554,g30216,g22125);
  or OR_16407(g30555,g30227,g22126);
  or OR_16408(g30556,g30236,g22127);
  or OR_16409(g30557,g30247,g22128);
  or OR_16410(g30558,g30258,g22129);
  or OR_16411(g30559,g30269,g22130);
  or OR_16412(g30560,g30278,g22131);
  or OR_16413(g30561,g30284,g22132);
  or OR_16414(g30562,g30289,g22133);
  or OR_16415(g30563,g29347,g22134);
  or OR_16416(g30579,g30173,g14571);
  or OR_16417(g30597,g13564,g29693);
  or OR_16418(g30605,g29529,g29520);
  or OR_16419(g30608,g13604,g29736);
  or OR_16420(g30609,g13633,g29742);
  or OR_16421(g30611,g13671,g29743);
  or OR_16422(g30672,g13737,g29752);
  or OR_16423(g30732,g13778,g29762);
  or OR_16424(g30733,g13807,g29773);
  or OR_16425(g30734,g13808,g29774);
  or OR_16426(g30824,g13833,g29789);
  or OR_16427(g30916,g13853,g29799);
  or OR_16428(g30984,g29765,g29755);
  or OR_16429(g31001,g29360,g28151);
  or OR_16430(g31002,g29362,g28154);
  or OR_16431(g31007,g29364,g28159);
  or OR_16432(g31014,g29367,g28160);
  or OR_16433(g31020,g29375,g28164);
  or OR_16434(g31144,g29477,g28193);
  or OR_16435(g31221,g29494,g28204);
  or OR_16436(g31241,g25959,g29510);
  or OR_16437(g31244,g25963,g29515);
  or OR_16438(g31245,g25964,g29516);
  or OR_16439(g31246,g25965,g29518);
  or OR_16440(g31247,g29513,g13324);
  or OR_16441(g31248,g25970,g29522);
  or OR_16442(g31249,g25971,g29523);
  or OR_16443(g31250,g25972,g29526);
  or OR_16444(g31251,g25973,g29527);
  or OR_16445(g31253,g25980,g29533);
  or OR_16446(g31254,g25981,g29534);
  or OR_16447(g31255,g25982,g29536);
  or OR_16448(g31256,g25983,g29537);
  or OR_16449(g31257,g29531,g28253);
  or OR_16450(g31258,g25991,g29550);
  or OR_16451(g31259,g25992,g29554);
  or OR_16452(g31260,g25993,g29555);
  or OR_16453(g31267,g29548,g28263);
  or OR_16454(g31268,g29552,g28266);
  or OR_16455(g31269,g26024,g29569);
  or OR_16456(g31274,g29565,g28280);
  or OR_16457(g31276,g29567,g28282);
  or OR_16458(g31277,g29570,g28285);
  or OR_16459(g31279,g29571,g29579);
  or OR_16460(g31284,g29575,g28290);
  or OR_16461(g31287,g29578,g28292);
  or OR_16462(g31288,g2955,g29914);
  or OR_16463(g31289,g29580,g29591);
  or OR_16464(g31291,g29581,g29593);
  or OR_16465(g31293,g29582,g28299);
  or OR_16466(g31295,g26090,g29598);
  or OR_16467(g31302,g29590,g28302);
  or OR_16468(g31303,g29592,g29606);
  or OR_16469(g31304,g29594,g29608);
  or OR_16470(g31306,g29595,g29610);
  or OR_16471(g31307,g29596,g28311);
  or OR_16472(g31308,g26101,g29614);
  or OR_16473(g31311,g26103,g29618);
  or OR_16474(g31315,g29607,g29623);
  or OR_16475(g31316,g29609,g29624);
  or OR_16476(g31317,g29611,g29626);
  or OR_16477(g31319,g29612,g28324);
  or OR_16478(g31320,g26125,g29632);
  or OR_16479(g31322,g26128,g29635);
  or OR_16480(g31325,g29625,g29639);
  or OR_16481(g31326,g29627,g29640);
  or OR_16482(g31375,g29628,g28339);
  or OR_16483(g31465,g26156,g29647);
  or OR_16484(g31466,g26160,g29650);
  or OR_16485(g31468,g29641,g29656);
  or OR_16486(g31472,g29642,g28352);
  or OR_16487(g31473,g26180,g29666);
  or OR_16488(g31474,g29668,g13583);
  or OR_16489(g31591,g29358,g29353);
  or OR_16490(g31668,g29924,g28558);
  or OR_16491(g31670,g29937,g28573);
  or OR_16492(g31745,g29959,g29973);
  or OR_16493(g31749,g29974,g29988);
  or OR_16494(g31751,g29975,g29990);
  or OR_16495(g31754,g29989,g30006);
  or OR_16496(g31755,g29991,g30008);
  or OR_16497(g31757,g29992,g30010);
  or OR_16498(g31760,g30007,g30027);
  or OR_16499(g31761,g30009,g30028);
  or OR_16500(g31762,g30011,g30030);
  or OR_16501(g31764,g30015,g30032);
  or OR_16502(g31766,g30029,g30042);
  or OR_16503(g31767,g30031,g30043);
  or OR_16504(g31768,g30033,g30045);
  or OR_16505(g31770,g30034,g30047);
  or OR_16506(g31772,g30035,g28654);
  or OR_16507(g31773,g30044,g30056);
  or OR_16508(g31774,g30046,g30057);
  or OR_16509(g31775,g30048,g30059);
  or OR_16510(g31779,g30050,g28673);
  or OR_16511(g31781,g30058,g30069);
  or OR_16512(g31782,g30060,g30070);
  or OR_16513(I29351,g29328,g29323,g29316,g30316);
  or OR_16514(I29352,g29322,g29315,g30315,g30308);
  or OR_16515(g31783,I29351,I29352);
  or OR_16516(g31785,g30071,g30082);
  or OR_16517(g31793,g28031,g30317);
  or OR_16518(g31864,g31271,g21703);
  or OR_16519(g31865,g31149,g21709);
  or OR_16520(g31866,g31252,g18142);
  or OR_16521(g31867,g31238,g18175);
  or OR_16522(g31868,g30600,g18204);
  or OR_16523(g31869,g30592,g18221);
  or OR_16524(g31870,g30607,g18262);
  or OR_16525(g31871,g30596,g18279);
  or OR_16526(g31872,g31524,g18535);
  or OR_16527(g31873,g31270,g21728);
  or OR_16528(g31874,g31016,g21729);
  or OR_16529(g31875,g31066,g21730);
  or OR_16530(g31876,g31125,g21731);
  or OR_16531(g31877,g31278,g21732);
  or OR_16532(g31878,g31015,g21733);
  or OR_16533(g31879,g31475,g21745);
  or OR_16534(g31880,g31280,g21774);
  or OR_16535(g31881,g31018,g21775);
  or OR_16536(g31882,g31115,g21776);
  or OR_16537(g31883,g31132,g21777);
  or OR_16538(g31884,g31290,g21778);
  or OR_16539(g31885,g31017,g21779);
  or OR_16540(g31886,g31481,g21791);
  or OR_16541(g31887,g31292,g21820);
  or OR_16542(g31888,g31067,g21821);
  or OR_16543(g31889,g31118,g21822);
  or OR_16544(g31890,g31143,g21823);
  or OR_16545(g31891,g31305,g21824);
  or OR_16546(g31892,g31019,g21825);
  or OR_16547(g31893,g31490,g21837);
  or OR_16548(g31894,g30671,g21870);
  or OR_16549(g31895,g31505,g24296);
  or OR_16550(g31896,g31242,g24305);
  or OR_16551(g31897,g31237,g24322);
  or OR_16552(g31898,g31707,g21906);
  or OR_16553(g31899,g31470,g21907);
  or OR_16554(g31900,g31484,g21908);
  or OR_16555(g31901,g31516,g21909);
  or OR_16556(g31902,g31744,g21910);
  or OR_16557(g31903,g31374,g21911);
  or OR_16558(g31904,g31780,g21923);
  or OR_16559(g31905,g31746,g21952);
  or OR_16560(g31906,g31477,g21953);
  or OR_16561(g31907,g31492,g21954);
  or OR_16562(g31908,g31519,g21955);
  or OR_16563(g31909,g31750,g21956);
  or OR_16564(g31910,g31471,g21957);
  or OR_16565(g31911,g31784,g21969);
  or OR_16566(g31912,g31752,g21998);
  or OR_16567(g31913,g31485,g21999);
  or OR_16568(g31914,g31499,g22000);
  or OR_16569(g31915,g31520,g22001);
  or OR_16570(g31916,g31756,g22002);
  or OR_16571(g31917,g31478,g22003);
  or OR_16572(g31918,g31786,g22015);
  or OR_16573(g31919,g31758,g22044);
  or OR_16574(g31920,g31493,g22045);
  or OR_16575(g31921,g31508,g22046);
  or OR_16576(g31922,g31525,g22047);
  or OR_16577(g31923,g31763,g22048);
  or OR_16578(g31924,g31486,g22049);
  or OR_16579(g31925,g31789,g22061);
  or OR_16580(g31926,g31765,g22090);
  or OR_16581(g31927,g31500,g22091);
  or OR_16582(g31928,g31517,g22092);
  or OR_16583(g31929,g31540,g22093);
  or OR_16584(g31930,g31769,g22094);
  or OR_16585(g31931,g31494,g22095);
  or OR_16586(g31932,g31792,g22107);
  or OR_16587(g31964,g31654,g14544);
  or OR_16588(g32037,g30566,g29329);
  or OR_16589(g32094,g30612,g29363);
  or OR_16590(g32117,g24482,g30914);
  or OR_16591(g32123,g30915,g30919);
  or OR_16592(g32124,g24488,g30920);
  or OR_16593(g32125,g30918,g29376);
  or OR_16594(g32130,g30921,g30925);
  or OR_16595(g32131,g24495,g30926);
  or OR_16596(g32132,g31487,g31479);
  or OR_16597(g32144,g30927,g30930);
  or OR_16598(g32155,g30935,g29475);
  or OR_16599(g32202,g31069,g13410);
  or OR_16600(g32208,g31120,g29584);
  or OR_16601(g32209,g31122,g29599);
  or OR_16602(g32210,g31123,g29600);
  or OR_16603(g32211,g31124,g29603);
  or OR_16604(g32216,g31128,g29615);
  or OR_16605(g32217,g31129,g29616);
  or OR_16606(g32218,g31130,g29619);
  or OR_16607(g32219,g31131,g29620);
  or OR_16608(g32220,g31139,g29633);
  or OR_16609(g32221,g31140,g29634);
  or OR_16610(g32222,g31141,g29636);
  or OR_16611(g32223,g31142,g29637);
  or OR_16612(g32225,g30576,g29336);
  or OR_16613(g32226,g31145,g29645);
  or OR_16614(g32227,g31146,g29648);
  or OR_16615(g32228,g31147,g29651);
  or OR_16616(g32229,g31148,g29652);
  or OR_16617(g32230,g30589,g29345);
  or OR_16618(g32231,g30590,g29346);
  or OR_16619(g32233,g31150,g29661);
  or OR_16620(g32235,g31151,g29662);
  or OR_16621(g32236,g31152,g29664);
  or OR_16622(g32237,g31153,g29667);
  or OR_16623(g32238,g30594,g29349);
  or OR_16624(g32239,g30595,g29350);
  or OR_16625(g32240,g24757,g31182);
  or OR_16626(g32243,g31166,g29683);
  or OR_16627(g32245,g31167,g29684);
  or OR_16628(g32247,g31168,g29686);
  or OR_16629(g32249,g31169,g29687);
  or OR_16630(g32250,g30598,g29351);
  or OR_16631(g32251,g30599,g29352);
  or OR_16632(g32252,g31183,g31206);
  or OR_16633(g32253,g24771,g31207);
  or OR_16634(g32257,g31184,g29708);
  or OR_16635(g32259,g31185,g29709);
  or OR_16636(g32262,g31186,g29710);
  or OR_16637(g32264,g31187,g29711);
  or OR_16638(g32266,g30604,g29354);
  or OR_16639(g32267,g31208,g31218);
  or OR_16640(g32268,g24785,g31219);
  or OR_16641(g32271,g31209,g29731);
  or OR_16642(g32275,g31210,g29732);
  or OR_16643(g32277,g31211,g29733);
  or OR_16644(g32279,g31220,g31224);
  or OR_16645(g32280,g24790,g31225);
  or OR_16646(g32285,g31222,g29740);
  or OR_16647(g32288,g31226,g31229);
  or OR_16648(g32289,g24796,g31230);
  or OR_16649(g32294,g31231,g31232);
  or OR_16650(g32344,g29804,g31266);
  or OR_16651(g32346,g29838,g31272);
  or OR_16652(g32347,g29839,g31273);
  or OR_16653(g32349,g29840,g31275);
  or OR_16654(g32351,g29851,g31281);
  or OR_16655(g32352,g29852,g31282);
  or OR_16656(g32353,g29853,g31283);
  or OR_16657(g32354,g29854,g31285);
  or OR_16658(g32355,g29855,g31286);
  or OR_16659(g32357,g29865,g31296);
  or OR_16660(g32358,g29866,g31297);
  or OR_16661(g32359,g29867,g31298);
  or OR_16662(g32360,g29868,g31299);
  or OR_16663(g32361,g29869,g31300);
  or OR_16664(g32362,g29870,g31301);
  or OR_16665(g32367,g29880,g31309);
  or OR_16666(g32368,g29881,g31310);
  or OR_16667(g32370,g29882,g31312);
  or OR_16668(g32371,g29883,g31313);
  or OR_16669(g32372,g29884,g31314);
  or OR_16670(g32373,g29894,g31321);
  or OR_16671(g32374,g29895,g31323);
  or OR_16672(g32375,g29896,g31324);
  or OR_16673(g32380,g29907,g31467);
  or OR_16674(g32385,g31480,g29938);
  or OR_16675(g32386,g31488,g29949);
  or OR_16676(g32387,g31489,g29952);
  or OR_16677(g32388,g31495,g29962);
  or OR_16678(g32389,g31496,g29966);
  or OR_16679(g32390,g31501,g29979);
  or OR_16680(g32391,g31502,g29982);
  or OR_16681(g32392,g31513,g30000);
  or OR_16682(g32395,g31523,g30049);
  or OR_16683(g32398,g31526,g30061);
  or OR_16684(g32399,g31527,g30062);
  or OR_16685(g32408,g31541,g30073);
  or OR_16686(g32426,g26105,g26131,g30613);
  or OR_16687(g32427,g8928,g30583);
  or OR_16688(g32429,g30318,g31794);
  or OR_16689(g32454,g30322,g31795);
  or OR_16690(I29985,g29385,g31376,g30735,g30825);
  or OR_16691(I29986,g31070,g31194,g30614,g30673);
  or OR_16692(I30054,g29385,g31376,g30735,g30825);
  or OR_16693(I30055,g31070,g31170,g30614,g30673);
  or OR_16694(I30123,g29385,g31376,g30735,g30825);
  or OR_16695(I30124,g31070,g31154,g30614,g30673);
  or OR_16696(I30192,g29385,g31376,g30735,g30825);
  or OR_16697(I30193,g31070,g30614,g30673,g31528);
  or OR_16698(I30261,g29385,g31376,g30735,g30825);
  or OR_16699(I30262,g31672,g31710,g31021,g30937);
  or OR_16700(I30330,g29385,g31376,g30735,g30825);
  or OR_16701(I30331,g31672,g31710,g31021,g30937);
  or OR_16702(I30399,g29385,g31376,g30735,g30825);
  or OR_16703(I30400,g31021,g30937,g31327,g30614);
  or OR_16704(I30468,g29385,g31376,g30735,g30825);
  or OR_16705(I30469,g31672,g31710,g31021,g30937);
  or OR_16706(g32976,g32207,g21704);
  or OR_16707(g32977,g32169,g21710);
  or OR_16708(g32978,g32197,g18145);
  or OR_16709(g32979,g32181,g18177);
  or OR_16710(g32980,g32254,g18198);
  or OR_16711(g32981,g32425,g18206);
  or OR_16712(g32982,g31948,g18208);
  or OR_16713(g32983,g31990,g18222);
  or OR_16714(g32984,g31934,g18264);
  or OR_16715(g32985,g31963,g18266);
  or OR_16716(g32986,g31996,g18280);
  or OR_16717(g32987,g32311,g18323);
  or OR_16718(g32988,g32232,g18325);
  or OR_16719(g32989,g32241,g18326);
  or OR_16720(g32990,g32281,g18341);
  or OR_16721(g32991,g32322,g18349);
  or OR_16722(g32992,g32242,g18351);
  or OR_16723(g32993,g32255,g18352);
  or OR_16724(g32994,g32290,g18367);
  or OR_16725(g32995,g32330,g18375);
  or OR_16726(g32996,g32256,g18377);
  or OR_16727(g32997,g32269,g18378);
  or OR_16728(g32998,g32300,g18393);
  or OR_16729(g32999,g32337,g18401);
  or OR_16730(g33000,g32270,g18403);
  or OR_16731(g33001,g32282,g18404);
  or OR_16732(g33002,g32304,g18419);
  or OR_16733(g33003,g32323,g18429);
  or OR_16734(g33004,g32246,g18431);
  or OR_16735(g33005,g32260,g18432);
  or OR_16736(g33006,g32291,g18447);
  or OR_16737(g33007,g32331,g18455);
  or OR_16738(g33008,g32261,g18457);
  or OR_16739(g33009,g32273,g18458);
  or OR_16740(g33010,g32301,g18473);
  or OR_16741(g33011,g32338,g18481);
  or OR_16742(g33012,g32274,g18483);
  or OR_16743(g33013,g32283,g18484);
  or OR_16744(g33014,g32305,g18499);
  or OR_16745(g33015,g32343,g18507);
  or OR_16746(g33016,g32284,g18509);
  or OR_16747(g33017,g32292,g18510);
  or OR_16748(g33018,g32312,g18525);
  or OR_16749(g33019,g32339,g18536);
  or OR_16750(g33020,g32160,g21734);
  or OR_16751(g33021,g32302,g21749);
  or OR_16752(g33022,g32306,g21750);
  or OR_16753(g33023,g32313,g21751);
  or OR_16754(g33024,g32324,g21752);
  or OR_16755(g33025,g32162,g21780);
  or OR_16756(g33026,g32307,g21795);
  or OR_16757(g33027,g32314,g21796);
  or OR_16758(g33028,g32325,g21797);
  or OR_16759(g33029,g32332,g21798);
  or OR_16760(g33030,g32166,g21826);
  or OR_16761(g33031,g32315,g21841);
  or OR_16762(g33032,g32326,g21842);
  or OR_16763(g33033,g32333,g21843);
  or OR_16764(g33034,g32340,g21844);
  or OR_16765(g33035,g32019,g21872);
  or OR_16766(g33036,g32168,g24309);
  or OR_16767(g33037,g32177,g24310);
  or OR_16768(g33038,g32184,g24311);
  or OR_16769(g33039,g32187,g24312);
  or OR_16770(g33040,g32164,g24313);
  or OR_16771(g33041,g32189,g24323);
  or OR_16772(g33042,g32193,g24324);
  or OR_16773(g33043,g32195,g24325);
  or OR_16774(g33044,g32199,g24327);
  or OR_16775(g33045,g32206,g24328);
  or OR_16776(g33046,g32308,g21912);
  or OR_16777(g33047,g31944,g21927);
  or OR_16778(g33048,g31960,g21928);
  or OR_16779(g33049,g31966,g21929);
  or OR_16780(g33050,g31974,g21930);
  or OR_16781(g33051,g32316,g21958);
  or OR_16782(g33052,g31961,g21973);
  or OR_16783(g33053,g31967,g21974);
  or OR_16784(g33054,g31975,g21975);
  or OR_16785(g33055,g31986,g21976);
  or OR_16786(g33056,g32327,g22004);
  or OR_16787(g33057,g31968,g22019);
  or OR_16788(g33058,g31976,g22020);
  or OR_16789(g33059,g31987,g22021);
  or OR_16790(g33060,g31992,g22022);
  or OR_16791(g33061,g32334,g22050);
  or OR_16792(g33062,g31977,g22065);
  or OR_16793(g33063,g31988,g22066);
  or OR_16794(g33064,g31993,g22067);
  or OR_16795(g33065,g32008,g22068);
  or OR_16796(g33066,g32341,g22096);
  or OR_16797(g33067,g31989,g22111);
  or OR_16798(g33068,g31994,g22112);
  or OR_16799(g33069,g32009,g22113);
  or OR_16800(g33070,g32010,g22114);
  or OR_16801(g33076,g32336,g32446);
  or OR_16802(g33115,g32397,g32401);
  or OR_16803(g33116,g32403,g32411);
  or OR_16804(g33118,g32413,g32418);
  or OR_16805(g33119,g32420,g32428);
  or OR_16806(g33123,g31962,g30577);
  or OR_16807(I30717,g31787,g32200,g31940,g31949);
  or OR_16808(I30718,g32348,g32356,g32097,g32020);
  or OR_16809(g33149,g32204,I30717,I30718);
  or OR_16810(g33159,g32016,g30730);
  or OR_16811(I30727,g31759,g32196,g31933,g31941);
  or OR_16812(I30728,g32345,g32350,g32056,g32018);
  or OR_16813(g33164,g32203,I30727,I30728);
  or OR_16814(I30734,g31790,g32191,g32086,g32095);
  or OR_16815(I30735,g32369,g32376,g32089,g32035);
  or OR_16816(g33176,g32198,I30734,I30735);
  or OR_16817(I30740,g31776,g32188,g32083,g32087);
  or OR_16818(I30741,g32085,g32030,g32224,g32013);
  or OR_16819(g33187,g32014,I30740,I30741);
  or OR_16820(I30745,g31777,g32321,g32069,g32084);
  or OR_16821(I30746,g32047,g31985,g31991,g32309);
  or OR_16822(g33197,g32342,I30745,I30746);
  or OR_16823(I30750,g31788,g32310,g32054,g32070);
  or OR_16824(I30751,g32042,g32161,g31943,g31959);
  or OR_16825(g33204,g32317,I30750,I30751);
  or OR_16826(I30755,g30564,g32303,g32049,g32055);
  or OR_16827(I30756,g32088,g32163,g32098,g32105);
  or OR_16828(g33212,g32328,I30755,I30756);
  or OR_16829(I30760,g31778,g32295,g32046,g32050);
  or OR_16830(I30761,g32071,g32167,g32067,g32082);
  or OR_16831(g33219,g32335,I30760,I30761);
  or OR_16832(g33227,g32029,g32031);
  or OR_16833(g33231,g32032,g32036);
  or OR_16834(g33232,g32034,g30936);
  or OR_16835(g33234,g32039,g32043);
  or OR_16836(g33235,g32040,g30982);
  or OR_16837(g33236,g32044,g32045);
  or OR_16838(g33238,g32048,g32051);
  or OR_16839(g33240,g32052,g32068);
  or OR_16840(g33251,g32096,g29509);
  or OR_16841(g33253,g32103,g29511);
  or OR_16842(g33254,g32104,g29512);
  or OR_16843(g33255,g32106,g29514);
  or OR_16844(g33256,g32107,g29517);
  or OR_16845(g33257,g32108,g29519);
  or OR_16846(g33259,g32109,g29521);
  or OR_16847(g33260,g32110,g29524);
  or OR_16848(g33261,g32111,g29525);
  or OR_16849(g33262,g32112,g29528);
  or OR_16850(g33265,g32113,g29530);
  or OR_16851(g33266,g32114,g29532);
  or OR_16852(g33267,g32115,g29535);
  or OR_16853(g33268,g32116,g29538);
  or OR_16854(g33270,g32119,g29547);
  or OR_16855(g33271,g32120,g29549);
  or OR_16856(g33272,g32121,g29551);
  or OR_16857(g33273,g32122,g29553);
  or OR_16858(g33274,g32126,g29563);
  or OR_16859(g33275,g32127,g29564);
  or OR_16860(g33276,g32128,g29566);
  or OR_16861(g33277,g32129,g29568);
  or OR_16862(g33278,g32139,g29572);
  or OR_16863(g33279,g32140,g29573);
  or OR_16864(g33280,g32141,g29574);
  or OR_16865(g33281,g32142,g29576);
  or OR_16866(g33282,g32143,g29577);
  or OR_16867(g33283,g31995,g30318);
  or OR_16868(g33286,g32145,g29585);
  or OR_16869(g33287,g32146,g29586);
  or OR_16870(g33288,g32147,g29587);
  or OR_16871(g33289,g32148,g29588);
  or OR_16872(g33290,g32149,g29589);
  or OR_16873(g33291,g32154,g13477);
  or OR_16874(g33292,g32150,g29601);
  or OR_16875(g33293,g32151,g29602);
  or OR_16876(g33294,g32152,g29604);
  or OR_16877(g33295,g32153,g29605);
  or OR_16878(g33296,g32156,g29617);
  or OR_16879(g33297,g32157,g29621);
  or OR_16880(g33298,g32158,g29622);
  or OR_16881(g33303,g32159,g29638);
  or OR_16882(g33310,g29631,g32165);
  or OR_16883(g33312,g29646,g32170);
  or OR_16884(g33313,g29649,g32171);
  or OR_16885(g33314,g29663,g32174);
  or OR_16886(g33315,g29665,g32175);
  or OR_16887(g33316,g29685,g32178);
  or OR_16888(g33317,g29688,g32179);
  or OR_16889(g33318,g31969,g32434);
  or OR_16890(g33321,g29712,g32182);
  or OR_16891(g33323,g31936,g32442);
  or OR_16892(g33380,g32234,g29926);
  or OR_16893(g33383,g32244,g29940);
  or OR_16894(g33384,g32248,g29943);
  or OR_16895(g33386,g32258,g29951);
  or OR_16896(g33387,g32263,g29954);
  or OR_16897(g33389,g32272,g29964);
  or OR_16898(g33390,g32276,g29968);
  or OR_16899(g33393,g32286,g29984);
  or OR_16900(g33534,g33186,g21700);
  or OR_16901(g33535,g33233,g21711);
  or OR_16902(g33536,g33241,g21715);
  or OR_16903(g33537,g33244,g21716);
  or OR_16904(g33538,g33252,g18144);
  or OR_16905(g33539,g33245,g18178);
  or OR_16906(g33540,g33099,g18207);
  or OR_16907(g33541,g33101,g18223);
  or OR_16908(g33542,g33102,g18265);
  or OR_16909(g33543,g33106,g18281);
  or OR_16910(g33544,g33392,g18317);
  or OR_16911(g33545,g33399,g18324);
  or OR_16912(g33546,g33402,g18327);
  or OR_16913(g33547,g33349,g18331);
  or OR_16914(g33548,g33327,g18336);
  or OR_16915(g33549,g33328,g18337);
  or OR_16916(g33550,g33342,g18338);
  or OR_16917(g33551,g33446,g18342);
  or OR_16918(g33552,g33400,g18343);
  or OR_16919(g33553,g33403,g18350);
  or OR_16920(g33554,g33407,g18353);
  or OR_16921(g33555,g33355,g18357);
  or OR_16922(g33556,g33329,g18362);
  or OR_16923(g33557,g33331,g18363);
  or OR_16924(g33558,g33350,g18364);
  or OR_16925(g33559,g33073,g18368);
  or OR_16926(g33560,g33404,g18369);
  or OR_16927(g33561,g33408,g18376);
  or OR_16928(g33562,g33414,g18379);
  or OR_16929(g33563,g33361,g18383);
  or OR_16930(g33564,g33332,g18388);
  or OR_16931(g33565,g33338,g18389);
  or OR_16932(g33566,g33356,g18390);
  or OR_16933(g33567,g33081,g18394);
  or OR_16934(g33568,g33409,g18395);
  or OR_16935(g33569,g33415,g18402);
  or OR_16936(g33570,g33420,g18405);
  or OR_16937(g33571,g33367,g18409);
  or OR_16938(g33572,g33339,g18414);
  or OR_16939(g33573,g33343,g18415);
  or OR_16940(g33574,g33362,g18416);
  or OR_16941(g33575,g33086,g18420);
  or OR_16942(g33576,g33401,g18423);
  or OR_16943(g33577,g33405,g18430);
  or OR_16944(g33578,g33410,g18433);
  or OR_16945(g33579,g33357,g18437);
  or OR_16946(g33580,g33330,g18442);
  or OR_16947(g33581,g33333,g18443);
  or OR_16948(g33582,g33351,g18444);
  or OR_16949(g33583,g33074,g18448);
  or OR_16950(g33584,g33406,g18449);
  or OR_16951(g33585,g33411,g18456);
  or OR_16952(g33586,g33416,g18459);
  or OR_16953(g33587,g33363,g18463);
  or OR_16954(g33588,g33334,g18468);
  or OR_16955(g33589,g33340,g18469);
  or OR_16956(g33590,g33358,g18470);
  or OR_16957(g33591,g33082,g18474);
  or OR_16958(g33592,g33412,g18475);
  or OR_16959(g33593,g33417,g18482);
  or OR_16960(g33594,g33421,g18485);
  or OR_16961(g33595,g33368,g18489);
  or OR_16962(g33596,g33341,g18494);
  or OR_16963(g33597,g33344,g18495);
  or OR_16964(g33598,g33364,g18496);
  or OR_16965(g33599,g33087,g18500);
  or OR_16966(g33600,g33418,g18501);
  or OR_16967(g33601,g33422,g18508);
  or OR_16968(g33602,g33425,g18511);
  or OR_16969(g33603,g33372,g18515);
  or OR_16970(g33604,g33345,g18520);
  or OR_16971(g33605,g33352,g18521);
  or OR_16972(g33606,g33369,g18522);
  or OR_16973(g33607,g33091,g18526);
  or OR_16974(g33608,g33322,g18537);
  or OR_16975(g33609,g33239,g18615);
  or OR_16976(g33610,g33242,g18616);
  or OR_16977(g33611,g33243,g18632);
  or OR_16978(g33612,g33247,g18633);
  or OR_16979(g33613,g33248,g18649);
  or OR_16980(g33614,g33249,g18650);
  or OR_16981(g33615,g33113,g21871);
  or OR_16982(g33616,g33237,g24314);
  or OR_16983(g33617,g33263,g24326);
  or OR_16984(g33618,g33353,g18757);
  or OR_16985(g33619,g33359,g18758);
  or OR_16986(g33620,g33360,g18774);
  or OR_16987(g33621,g33365,g18775);
  or OR_16988(g33622,g33366,g18791);
  or OR_16989(g33623,g33370,g18792);
  or OR_16990(g33624,g33371,g18808);
  or OR_16991(g33625,g33373,g18809);
  or OR_16992(g33626,g33374,g18825);
  or OR_16993(g33627,g33376,g18826);
  or OR_16994(g33628,g33071,g32450);
  or OR_16995(g33685,g32396,g33423);
  or OR_16996(g33692,g32400,g33428);
  or OR_16997(g33694,g32402,g33429);
  or OR_16998(g33699,g32409,g33433);
  or OR_16999(g33703,g32410,g33434);
  or OR_17000(g33706,g32412,g33440);
  or OR_17001(g33709,g32414,g33441);
  or OR_17002(g33714,g32419,g33450);
  or OR_17003(g33732,g33104,g32011);
  or OR_17004(g33733,g33105,g32012);
  or OR_17005(g33788,g33122,g32041);
  or OR_17006(g33791,g33379,g32430);
  or OR_17007(g33794,g33126,g32053);
  or OR_17008(g33891,g33264,g33269);
  or OR_17009(g33914,g33305,g33311);
  or OR_17010(g33945,g32430,g33455);
  or OR_17011(g33946,g32434,g33456);
  or OR_17012(g33947,g32438,g33457);
  or OR_17013(g33948,g32442,g33458);
  or OR_17014(g33949,g32446,g33459);
  or OR_17015(g33950,g32450,g33460);
  or OR_17016(I31838,g33461,g33462,g33463,g33464);
  or OR_17017(I31839,g33465,g33466,g33467,g33468);
  or OR_17018(g33951,g33469,I31838,I31839);
  or OR_17019(I31843,g33470,g33471,g33472,g33473);
  or OR_17020(I31844,g33474,g33475,g33476,g33477);
  or OR_17021(g33952,g33478,I31843,I31844);
  or OR_17022(I31848,g33479,g33480,g33481,g33482);
  or OR_17023(I31849,g33483,g33484,g33485,g33486);
  or OR_17024(g33953,g33487,I31848,I31849);
  or OR_17025(I31853,g33488,g33489,g33490,g33491);
  or OR_17026(I31854,g33492,g33493,g33494,g33495);
  or OR_17027(g33954,g33496,I31853,I31854);
  or OR_17028(I31858,g33497,g33498,g33499,g33500);
  or OR_17029(I31859,g33501,g33502,g33503,g33504);
  or OR_17030(g33955,g33505,I31858,I31859);
  or OR_17031(I31863,g33506,g33507,g33508,g33509);
  or OR_17032(I31864,g33510,g33511,g33512,g33513);
  or OR_17033(g33956,g33514,I31863,I31864);
  or OR_17034(I31868,g33515,g33516,g33517,g33518);
  or OR_17035(I31869,g33519,g33520,g33521,g33522);
  or OR_17036(g33957,g33523,I31868,I31869);
  or OR_17037(I31873,g33524,g33525,g33526,g33527);
  or OR_17038(I31874,g33528,g33529,g33530,g33531);
  or OR_17039(g33958,g33532,I31873,I31874);
  or OR_17040(g33960,g33759,g21701);
  or OR_17041(g33961,g33789,g21712);
  or OR_17042(g33962,g33822,g18123);
  or OR_17043(g33963,g33830,g18124);
  or OR_17044(g33964,g33817,g18146);
  or OR_17045(g33965,g33805,g18179);
  or OR_17046(g33966,g33837,g18318);
  or OR_17047(g33967,g33842,g18319);
  or OR_17048(g33968,g33855,g18320);
  or OR_17049(g33969,g33864,g18321);
  or OR_17050(g33970,g33868,g18322);
  or OR_17051(g33971,g33890,g18330);
  or OR_17052(g33972,g33941,g18335);
  or OR_17053(g33973,g33840,g18344);
  or OR_17054(g33974,g33846,g18345);
  or OR_17055(g33975,g33860,g18346);
  or OR_17056(g33976,g33869,g18347);
  or OR_17057(g33977,g33876,g18348);
  or OR_17058(g33978,g33892,g18356);
  or OR_17059(g33979,g33942,g18361);
  or OR_17060(g33980,g33843,g18370);
  or OR_17061(g33981,g33856,g18371);
  or OR_17062(g33982,g33865,g18372);
  or OR_17063(g33983,g33877,g18373);
  or OR_17064(g33984,g33881,g18374);
  or OR_17065(g33985,g33896,g18382);
  or OR_17066(g33986,g33639,g18387);
  or OR_17067(g33987,g33847,g18396);
  or OR_17068(g33988,g33861,g18397);
  or OR_17069(g33989,g33870,g18398);
  or OR_17070(g33990,g33882,g18399);
  or OR_17071(g33991,g33885,g18400);
  or OR_17072(g33992,g33900,g18408);
  or OR_17073(g33993,g33646,g18413);
  or OR_17074(g33994,g33841,g18424);
  or OR_17075(g33995,g33848,g18425);
  or OR_17076(g33996,g33862,g18426);
  or OR_17077(g33997,g33871,g18427);
  or OR_17078(g33998,g33878,g18428);
  or OR_17079(g33999,g33893,g18436);
  or OR_17080(g34000,g33943,g18441);
  or OR_17081(g34001,g33844,g18450);
  or OR_17082(g34002,g33857,g18451);
  or OR_17083(g34003,g33866,g18452);
  or OR_17084(g34004,g33879,g18453);
  or OR_17085(g34005,g33883,g18454);
  or OR_17086(g34006,g33897,g18462);
  or OR_17087(g34007,g33640,g18467);
  or OR_17088(g34008,g33849,g18476);
  or OR_17089(g34009,g33863,g18477);
  or OR_17090(g34010,g33872,g18478);
  or OR_17091(g34011,g33884,g18479);
  or OR_17092(g34012,g33886,g18480);
  or OR_17093(g34013,g33901,g18488);
  or OR_17094(g34014,g33647,g18493);
  or OR_17095(g34015,g33858,g18502);
  or OR_17096(g34016,g33867,g18503);
  or OR_17097(g34017,g33880,g18504);
  or OR_17098(g34018,g33887,g18505);
  or OR_17099(g34019,g33889,g18506);
  or OR_17100(g34020,g33904,g18514);
  or OR_17101(g34021,g33652,g18519);
  or OR_17102(g34022,g33873,g18538);
  or OR_17103(g34023,g33796,g24320);
  or OR_17104(g34024,g33807,g24331);
  or OR_17105(g34025,g33927,g18672);
  or OR_17106(g34026,g33715,g18682);
  or OR_17107(g34027,g33718,g18683);
  or OR_17108(g34028,g33720,g18684);
  or OR_17109(g34029,g33798,g18703);
  or OR_17110(g34030,g33727,g18704);
  or OR_17111(g34031,g33735,g18705);
  or OR_17112(g34032,g33816,g18706);
  or OR_17113(g34033,g33821,g18708);
  or OR_17114(g34034,g33719,g18713);
  or OR_17115(g34035,g33721,g18714);
  or OR_17116(g34036,g33722,g18715);
  or OR_17117(g34037,g33803,g18734);
  or OR_17118(g34038,g33731,g18735);
  or OR_17119(g34039,g33743,g18736);
  or OR_17120(g34040,g33818,g18737);
  or OR_17121(g34041,g33829,g18739);
  or OR_17122(g34043,g33903,g33905);
  or OR_17123(g34046,g33906,g33908);
  or OR_17124(g34055,g33909,g33910);
  or OR_17125(g34057,g33911,g33915);
  or OR_17126(g34064,g33919,g33922);
  or OR_17127(g34090,g33676,g33680);
  or OR_17128(g34095,g33681,g33687);
  or OR_17129(g34099,g33684,g33689);
  or OR_17130(g34100,g33690,g33697);
  or OR_17131(g34101,g33693,g33700);
  or OR_17132(g34103,g33701,g33707);
  or OR_17133(g34107,g33710,g33121);
  or OR_17134(g34125,g33724,g33124);
  or OR_17135(g34127,g33657,g32438);
  or OR_17136(g34148,g33758,g19656);
  or OR_17137(g34149,g33760,g19674);
  or OR_17138(g34153,g33899,g33451);
  or OR_17139(g34158,g33784,g19740);
  or OR_17140(g34166,g33785,g19752);
  or OR_17141(g34167,g33786,g19768);
  or OR_17142(g34168,g33787,g19784);
  or OR_17143(g34170,g33790,g19855);
  or OR_17144(g34172,g33795,g19914);
  or OR_17145(g34189,g33801,g33808);
  or OR_17146(g34190,g33802,g33810);
  or OR_17147(g34193,g33809,g33814);
  or OR_17148(g34194,g33811,g33815);
  or OR_17149(g34199,g33820,g33828);
  or OR_17150(g34204,g33832,g33833);
  or OR_17151(g34206,g33834,g33836);
  or OR_17152(g34207,g33835,g33304);
  or OR_17153(g34231,g33898,g33902);
  or OR_17154(g34232,g33451,g33944);
  or OR_17155(g34233,g32455,g33951);
  or OR_17156(g34234,g32520,g33952);
  or OR_17157(g34235,g32585,g33953);
  or OR_17158(g34236,g32650,g33954);
  or OR_17159(g34237,g32715,g33955);
  or OR_17160(g34238,g32780,g33956);
  or OR_17161(g34239,g32845,g33957);
  or OR_17162(g34240,g32910,g33958);
  or OR_17163(g34249,g34110,g21702);
  or OR_17164(g34250,g34111,g21713);
  or OR_17165(g34251,g34157,g18147);
  or OR_17166(g34252,g34146,g18180);
  or OR_17167(g34253,g34171,g24300);
  or OR_17168(g34254,g34116,g24301);
  or OR_17169(g34255,g34120,g24302);
  or OR_17170(g34256,g34173,g24303);
  or OR_17171(g34257,g34226,g18674);
  or OR_17172(g34258,g34211,g18675);
  or OR_17173(g34259,g34066,g18679);
  or OR_17174(g34260,g34113,g18680);
  or OR_17175(g34261,g34074,g18688);
  or OR_17176(g34262,g34075,g18697);
  or OR_17177(g34263,g34078,g18699);
  or OR_17178(g34264,g34081,g18701);
  or OR_17179(g34265,g34117,g18711);
  or OR_17180(g34266,g34076,g18719);
  or OR_17181(g34267,g34079,g18728);
  or OR_17182(g34268,g34082,g18730);
  or OR_17183(g34269,g34083,g18732);
  or OR_17184(g34273,g27765,g34203);
  or OR_17185(g34274,g27822,g34205);
  or OR_17186(g34278,g26829,g34212);
  or OR_17187(g34280,g26833,g34213);
  or OR_17188(g34282,g26838,g34214);
  or OR_17189(g34283,g26839,g34215);
  or OR_17190(g34286,g26842,g34216);
  or OR_17191(g34288,g26846,g34217);
  or OR_17192(g34289,g26847,g34218);
  or OR_17193(g34290,g26848,g34219);
  or OR_17194(g34292,g26853,g34223);
  or OR_17195(g34293,g26854,g34224);
  or OR_17196(g34294,g26855,g34225);
  or OR_17197(g34297,g26858,g34228);
  or OR_17198(g34300,g26864,g34230);
  or OR_17199(g34303,g25768,g34045);
  or OR_17200(g34305,g25775,g34050);
  or OR_17201(g34306,g25782,g34054);
  or OR_17202(g34314,g25831,g34061);
  or OR_17203(g34318,g25850,g34063);
  or OR_17204(g34321,g25866,g34065);
  or OR_17205(g34330,g34069,g33717);
  or OR_17206(g34331,g27121,g34072);
  or OR_17207(g34332,g34071,g33723);
  or OR_17208(g34347,g25986,g34102);
  or OR_17209(g34349,g26019,g34104);
  or OR_17210(g34350,g26048,g34106);
  or OR_17211(g34352,g26079,g34109);
  or OR_17212(g34353,g26088,g34114);
  or OR_17213(g34366,g26257,g34133);
  or OR_17214(g34368,g26274,g34135);
  or OR_17215(g34369,g26279,g34136);
  or OR_17216(g34372,g26287,g34137);
  or OR_17217(g34373,g26292,g34138);
  or OR_17218(g34374,g26294,g34139);
  or OR_17219(g34376,g26301,g34140);
  or OR_17220(g34377,g26304,g34141);
  or OR_17221(g34379,g26312,g34143);
  or OR_17222(g34399,g34178,g25067);
  or OR_17223(g34402,g34179,g25084);
  or OR_17224(g34403,g34180,g25085);
  or OR_17225(g34404,g34182,g25102);
  or OR_17226(g34405,g34183,g25103);
  or OR_17227(g34406,g34184,g25123);
  or OR_17228(g34407,g34185,g25124);
  or OR_17229(g34411,g34186,g25142);
  or OR_17230(g34412,g34187,g25143);
  or OR_17231(g34416,g34191,g25159);
  or OR_17232(g34417,g27678,g34196);
  or OR_17233(g34421,g27686,g34198);
  or OR_17234(g34438,g34348,g18150);
  or OR_17235(g34439,g34344,g18181);
  or OR_17236(g34440,g34364,g24226);
  or OR_17237(g34441,g34381,g18540);
  or OR_17238(g34442,g34380,g18542);
  or OR_17239(g34443,g34385,g18545);
  or OR_17240(g34444,g34389,g18546);
  or OR_17241(g34445,g34382,g18548);
  or OR_17242(g34446,g34390,g18550);
  or OR_17243(g34447,g34363,g18552);
  or OR_17244(g34448,g34365,g18553);
  or OR_17245(g34449,g34279,g18662);
  or OR_17246(g34450,g34281,g18663);
  or OR_17247(g34451,g34393,g18664);
  or OR_17248(g34452,g34401,g18665);
  or OR_17249(g34453,g34410,g18666);
  or OR_17250(g34454,g34414,g18667);
  or OR_17251(g34455,g34284,g18668);
  or OR_17252(g34456,g34395,g18669);
  or OR_17253(g34457,g34394,g18670);
  or OR_17254(g34458,g34396,g18671);
  or OR_17255(g34459,g34415,g18673);
  or OR_17256(g34460,g34301,g18677);
  or OR_17257(g34461,g34291,g18681);
  or OR_17258(g34462,g34334,g18685);
  or OR_17259(g34463,g34338,g18686);
  or OR_17260(g34464,g34340,g18687);
  or OR_17261(g34465,g34295,g18712);
  or OR_17262(g34466,g34337,g18716);
  or OR_17263(g34467,g34341,g18717);
  or OR_17264(g34468,g34342,g18718);
  or OR_17265(g34494,g26849,g34413);
  or OR_17266(g34535,g34309,g34073);
  or OR_17267(g34537,g34324,g34084);
  or OR_17268(g34598,g34541,g18136);
  or OR_17269(g34599,g34542,g18149);
  or OR_17270(g34600,g34538,g18182);
  or OR_17271(g34601,g34488,g18211);
  or OR_17272(g34602,g34489,g18269);
  or OR_17273(g34603,g34561,g15075);
  or OR_17274(g34604,g34563,g15076);
  or OR_17275(g34605,g34566,g15077);
  or OR_17276(g34606,g34564,g15080);
  or OR_17277(g34607,g34567,g15081);
  or OR_17278(g34608,g34568,g15082);
  or OR_17279(g34609,g34503,g18563);
  or OR_17280(g34610,g34507,g18564);
  or OR_17281(g34611,g34508,g18565);
  or OR_17282(g34612,g34514,g18566);
  or OR_17283(g34613,g34515,g18567);
  or OR_17284(g34614,g34518,g18568);
  or OR_17285(g34615,g34516,g18576);
  or OR_17286(g34616,g34519,g18577);
  or OR_17287(g34617,g34526,g18579);
  or OR_17288(g34618,g34527,g18580);
  or OR_17289(g34619,g34528,g18581);
  or OR_17290(g34620,g34529,g18582);
  or OR_17291(g34621,g34517,g18583);
  or OR_17292(g34622,g34520,g18584);
  or OR_17293(g34623,g34525,g18585);
  or OR_17294(g34624,g34509,g18592);
  or OR_17295(g34625,g34532,g18610);
  or OR_17296(g34626,g34533,g18627);
  or OR_17297(g34627,g34534,g18644);
  or OR_17298(g34628,g34493,g18653);
  or OR_17299(g34629,g34495,g18654);
  or OR_17300(g34630,g34560,g15117);
  or OR_17301(g34631,g34562,g15118);
  or OR_17302(g34632,g34565,g15119);
  or OR_17303(g34633,g34481,g18690);
  or OR_17304(g34634,g34483,g18691);
  or OR_17305(g34635,g34485,g18692);
  or OR_17306(g34636,g34476,g18693);
  or OR_17307(g34637,g34478,g18694);
  or OR_17308(g34638,g34484,g18721);
  or OR_17309(g34639,g34486,g18722);
  or OR_17310(g34640,g34487,g18723);
  or OR_17311(g34641,g34479,g18724);
  or OR_17312(g34642,g34482,g18725);
  or OR_17313(g34643,g34554,g18752);
  or OR_17314(g34644,g34555,g18769);
  or OR_17315(g34645,g34556,g18786);
  or OR_17316(g34646,g34557,g18803);
  or OR_17317(g34647,g34558,g18820);
  or OR_17318(g34649,g33111,g34492);
  or OR_17319(g34657,g33114,g34497);
  or OR_17320(g34663,g32028,g34500);
  or OR_17321(g34693,g34513,g34310);
  or OR_17322(g34695,g34523,g34322);
  or OR_17323(g34708,g33381,g34572);
  or OR_17324(g34719,g34701,g18133);
  or OR_17325(g34720,g34694,g18134);
  or OR_17326(g34721,g34696,g18135);
  or OR_17327(g34722,g34707,g18137);
  or OR_17328(g34723,g34710,g18139);
  or OR_17329(g34724,g34702,g18152);
  or OR_17330(g34725,g34700,g18183);
  or OR_17331(g34726,g34665,g18212);
  or OR_17332(g34727,g34655,g18213);
  or OR_17333(g34728,g34661,g18214);
  or OR_17334(g34729,g34666,g18270);
  or OR_17335(g34730,g34658,g18271);
  or OR_17336(g34731,g34662,g18272);
  or OR_17337(g34732,g34686,g18593);
  or OR_17338(g34733,g34678,g18651);
  or OR_17339(g34734,g34681,g18652);
  or OR_17340(g34735,g34709,g15116);
  or OR_17341(g34761,g34679,g34506);
  or OR_17342(g34762,g34687,g34524);
  or OR_17343(g34781,g33431,g34715);
  or OR_17344(g34783,g33110,g34667);
  or OR_17345(g34790,g34774,g18151);
  or OR_17346(g34791,g34771,g18184);
  or OR_17347(g34792,g34750,g18569);
  or OR_17348(g34793,g34744,g18570);
  or OR_17349(g34794,g34746,g18571);
  or OR_17350(g34795,g34753,g18572);
  or OR_17351(g34796,g34745,g18573);
  or OR_17352(g34797,g34747,g18574);
  or OR_17353(g34798,g34754,g18575);
  or OR_17354(g34799,g34751,g18578);
  or OR_17355(g34800,g34752,g18586);
  or OR_17356(g34801,g34756,g18588);
  or OR_17357(g34802,g34757,g18589);
  or OR_17358(g34803,g34758,g18590);
  or OR_17359(g34804,g34740,g18591);
  or OR_17360(g34805,g34748,g18594);
  or OR_17361(g34806,g34763,g18595);
  or OR_17362(g34807,g34764,g18596);
  or OR_17363(g34808,g34765,g18599);
  or OR_17364(g34809,g33677,g34738);
  or OR_17365(g34819,g34741,g34684);
  or OR_17366(g34826,g34742,g34685);
  or OR_17367(g34843,g33924,g34782);
  or OR_17368(g34849,g34842,g18154);
  or OR_17369(g34850,g34841,g18185);
  or OR_17370(g34856,g34811,g34743);
  or OR_17371(g34880,g34867,g18153);
  or OR_17372(g34881,g34866,g18187);
  or OR_17373(g34882,g34876,g18659);
  or OR_17374(g34884,g34858,g21666);
  or OR_17375(g34887,g34865,g21670);
  or OR_17376(g34890,g34863,g21674);
  or OR_17377(g34894,g34862,g21678);
  or OR_17378(g34897,g34861,g21682);
  or OR_17379(g34900,g34860,g21686);
  or OR_17380(g34903,g34859,g21690);
  or OR_17381(g34906,g34857,g21694);
  or OR_17382(g34911,g34909,g18188);
  or OR_17383(g34931,g2984,g34912);
  or OR_17384(g34957,g34948,g21662);
  or OR_17385(g34970,g34868,g34961);
  or OR_17386(g34971,g34869,g34962);
  or OR_17387(g34974,g34870,g34963);
  or OR_17388(g34975,g34871,g34964);
  or OR_17389(g34976,g34872,g34965);
  or OR_17390(g34977,g34873,g34966);
  or OR_17391(g34978,g34874,g34967);
  or OR_17392(g34979,g34875,g34968);
  or OR_17393(g34980,g34969,g18587);
  or OR_17394(g35000,g34953,g34999);
  nand NAND_17395(I11824,g4593,g4601);
  nand NAND_17396(I11825,g4593,I11824);
  nand NAND_17397(I11826,g4601,I11824);
  nand NAND_17398(g7133,I11825,I11826);
  nand NAND_17399(g7150,g5016,g5062);
  nand NAND_17400(g7167,g5360,g5406);
  nand NAND_17401(g7184,g5706,g5752);
  nand NAND_17402(I11864,g4434,g4401);
  nand NAND_17403(I11865,g4434,I11864);
  nand NAND_17404(I11866,g4401,I11864);
  nand NAND_17405(g7201,I11865,I11866);
  nand NAND_17406(g7209,g6052,g6098);
  nand NAND_17407(I11877,g4388,g4430);
  nand NAND_17408(I11878,g4388,I11877);
  nand NAND_17409(I11879,g4430,I11877);
  nand NAND_17410(g7223,I11878,I11879);
  nand NAND_17411(g7227,g4584,g4593);
  nand NAND_17412(g7228,g6398,g6444);
  nand NAND_17413(g7442,g896,g890);
  nand NAND_17414(g7549,g1018,g1030);
  nand NAND_17415(g7582,g1361,g1373);
  nand NAND_17416(I12074,g996,g979);
  nand NAND_17417(I12075,g996,I12074);
  nand NAND_17418(I12076,g979,I12074);
  nand NAND_17419(g7598,I12075,I12076);
  nand NAND_17420(g7611,g4057,g4064);
  nand NAND_17421(I12096,g1339,g1322);
  nand NAND_17422(I12097,g1339,I12096);
  nand NAND_17423(I12098,g1322,I12096);
  nand NAND_17424(g7620,I12097,I12098);
  nand NAND_17425(g7690,g4669,g4659,g4653);
  nand NAND_17426(g7701,g4859,g4849,g4843);
  nand NAND_17427(I12203,g1094,g1135);
  nand NAND_17428(I12204,g1094,I12203);
  nand NAND_17429(I12205,g1135,I12203);
  nand NAND_17430(g7803,I12204,I12205);
  nand NAND_17431(I12217,g1437,g1478);
  nand NAND_17432(I12218,g1437,I12217);
  nand NAND_17433(I12219,g1478,I12217);
  nand NAND_17434(g7823,I12218,I12219);
  nand NAND_17435(g7836,g4653,g4688);
  nand NAND_17436(g7846,g4843,g4878);
  nand NAND_17437(g7850,g554,g807);
  nand NAND_17438(I12240,g1111,g1105);
  nand NAND_17439(I12241,g1111,I12240);
  nand NAND_17440(I12242,g1105,I12240);
  nand NAND_17441(g7857,I12241,I12242);
  nand NAND_17442(I12251,g1124,g1129);
  nand NAND_17443(I12252,g1124,I12251);
  nand NAND_17444(I12253,g1129,I12251);
  nand NAND_17445(g7869,I12252,I12253);
  nand NAND_17446(I12261,g1454,g1448);
  nand NAND_17447(I12262,g1454,I12261);
  nand NAND_17448(I12263,g1448,I12261);
  nand NAND_17449(g7879,I12262,I12263);
  nand NAND_17450(I12269,g1141,g956);
  nand NAND_17451(I12270,g1141,I12269);
  nand NAND_17452(I12271,g956,I12269);
  nand NAND_17453(g7885,I12270,I12271);
  nand NAND_17454(I12277,g1467,g1472);
  nand NAND_17455(I12278,g1467,I12277);
  nand NAND_17456(I12279,g1472,I12277);
  nand NAND_17457(g7887,I12278,I12279);
  nand NAND_17458(I12287,g1484,g1300);
  nand NAND_17459(I12288,g1484,I12287);
  nand NAND_17460(I12289,g1300,I12287);
  nand NAND_17461(g7897,I12288,I12289);
  nand NAND_17462(I12344,g3106,g3111);
  nand NAND_17463(I12345,g3106,I12344);
  nand NAND_17464(I12346,g3111,I12344);
  nand NAND_17465(g8010,I12345,I12346);
  nand NAND_17466(I12372,g3457,g3462);
  nand NAND_17467(I12373,g3457,I12372);
  nand NAND_17468(I12374,g3462,I12372);
  nand NAND_17469(g8069,I12373,I12374);
  nand NAND_17470(g8105,g3068,g3072);
  nand NAND_17471(I12401,g3808,g3813);
  nand NAND_17472(I12402,g3808,I12401);
  nand NAND_17473(I12403,g3813,I12401);
  nand NAND_17474(g8124,I12402,I12403);
  nand NAND_17475(g8163,g3419,g3423);
  nand NAND_17476(g8227,g3770,g3774);
  nand NAND_17477(I12468,g405,g392);
  nand NAND_17478(I12469,g405,I12468);
  nand NAND_17479(I12470,g392,I12468);
  nand NAND_17480(g8238,I12469,I12470);
  nand NAND_17481(g8292,g218,g215);
  nand NAND_17482(g8347,g4358,g4349,g4340);
  nand NAND_17483(I12544,g191,g194);
  nand NAND_17484(I12545,g191,I12544);
  nand NAND_17485(I12546,g194,I12544);
  nand NAND_17486(g8359,I12545,I12546);
  nand NAND_17487(g8434,g3080,g3072);
  nand NAND_17488(g8500,g3431,g3423);
  nand NAND_17489(g8561,g3782,g3774);
  nand NAND_17490(g8609,g1171,g1157);
  nand NAND_17491(g8632,g1514,g1500);
  nand NAND_17492(g8678,g376,g358);
  nand NAND_17493(g8691,g3267,g3310,g3281,g3303);
  nand NAND_17494(g8728,g3618,g3661,g3632,g3654);
  nand NAND_17495(I12728,g4291,g4287);
  nand NAND_17496(I12729,g4291,I12728);
  nand NAND_17497(I12730,g4287,I12728);
  nand NAND_17498(g8737,I12729,I12730);
  nand NAND_17499(g8751,g3969,g4012,g3983,g4005);
  nand NAND_17500(g8769,g691,g714);
  nand NAND_17501(g8803,g128,g4646);
  nand NAND_17502(g8806,g358,g370,g376,g385);
  nand NAND_17503(g8829,g5011,g4836);
  nand NAND_17504(g8847,g4831,g4681);
  nand NAND_17505(I12840,g4222,g4235);
  nand NAND_17506(I12841,g4222,I12840);
  nand NAND_17507(I12842,g4235,I12840);
  nand NAND_17508(g8871,I12841,I12842);
  nand NAND_17509(I12848,g4281,g4277);
  nand NAND_17510(I12849,g4281,I12848);
  nand NAND_17511(I12850,g4277,I12848);
  nand NAND_17512(g8873,I12849,I12850);
  nand NAND_17513(g8889,g3684,g4871);
  nand NAND_17514(I12876,g4200,g4180);
  nand NAND_17515(I12877,g4200,I12876);
  nand NAND_17516(I12878,g4180,I12876);
  nand NAND_17517(g8913,I12877,I12878);
  nand NAND_17518(g8967,g4264,g4258);
  nand NAND_17519(g9092,g3004,g3050);
  nand NAND_17520(g9177,g3355,g3401);
  nand NAND_17521(g9203,g3706,g3752);
  nand NAND_17522(g9246,g847,g812);
  nand NAND_17523(I13043,g5115,g5120);
  nand NAND_17524(I13044,g5115,I13043);
  nand NAND_17525(I13045,g5120,I13043);
  nand NAND_17526(g9258,I13044,I13045);
  nand NAND_17527(I13065,g4308,g4304);
  nand NAND_17528(I13066,g4308,I13065);
  nand NAND_17529(I13067,g4304,I13065);
  nand NAND_17530(g9295,I13066,I13067);
  nand NAND_17531(I13077,g5462,g5467);
  nand NAND_17532(I13078,g5462,I13077);
  nand NAND_17533(I13079,g5467,I13077);
  nand NAND_17534(g9310,I13078,I13079);
  nand NAND_17535(g9334,g827,g832);
  nand NAND_17536(g9372,g5080,g5084);
  nand NAND_17537(I13109,g5808,g5813);
  nand NAND_17538(I13110,g5808,I13109);
  nand NAND_17539(I13111,g5813,I13109);
  nand NAND_17540(g9391,I13110,I13111);
  nand NAND_17541(g9442,g5424,g5428);
  nand NAND_17542(I13139,g6154,g6159);
  nand NAND_17543(I13140,g6154,I13139);
  nand NAND_17544(I13141,g6159,I13139);
  nand NAND_17545(g9461,I13140,I13141);
  nand NAND_17546(g9485,g1657,g1624);
  nand NAND_17547(g9509,g5770,g5774);
  nand NAND_17548(I13182,g6500,g6505);
  nand NAND_17549(I13183,g6500,I13182);
  nand NAND_17550(I13184,g6505,I13182);
  nand NAND_17551(g9528,I13183,I13184);
  nand NAND_17552(g9538,g1792,g1760);
  nand NAND_17553(g9543,g2217,g2185);
  nand NAND_17554(g9567,g6116,g6120);
  nand NAND_17555(g9591,g1926,g1894);
  nand NAND_17556(g9595,g2351,g2319);
  nand NAND_17557(g9629,g6462,g6466);
  nand NAND_17558(g9645,g2060,g2028);
  nand NAND_17559(g9654,g2485,g2453);
  nand NAND_17560(g9663,g128,g4646);
  nand NAND_17561(g9705,g2619,g2587);
  nand NAND_17562(g9715,g5011,g4836);
  nand NAND_17563(g9724,g5092,g5084);
  nand NAND_17564(I13334,g1687,g1691);
  nand NAND_17565(I13335,g1687,I13334);
  nand NAND_17566(I13336,g1691,I13334);
  nand NAND_17567(g9750,I13335,I13336);
  nand NAND_17568(g9775,g4831,g4681);
  nand NAND_17569(g9800,g5436,g5428);
  nand NAND_17570(I13382,g269,g246);
  nand NAND_17571(I13383,g269,I13382);
  nand NAND_17572(I13384,g246,I13382);
  nand NAND_17573(g9823,I13383,I13384);
  nand NAND_17574(I13390,g1821,g1825);
  nand NAND_17575(I13391,g1821,I13390);
  nand NAND_17576(I13392,g1825,I13390);
  nand NAND_17577(g9825,I13391,I13392);
  nand NAND_17578(I13401,g2246,g2250);
  nand NAND_17579(I13402,g2246,I13401);
  nand NAND_17580(I13403,g2250,I13401);
  nand NAND_17581(g9830,I13402,I13403);
  nand NAND_17582(g9852,g3684,g4871);
  nand NAND_17583(g9883,g5782,g5774);
  nand NAND_17584(I13442,g262,g239);
  nand NAND_17585(I13443,g262,I13442);
  nand NAND_17586(I13444,g239,I13442);
  nand NAND_17587(g9904,I13443,I13444);
  nand NAND_17588(I13452,g1955,g1959);
  nand NAND_17589(I13453,g1955,I13452);
  nand NAND_17590(I13454,g1959,I13452);
  nand NAND_17591(g9908,I13453,I13454);
  nand NAND_17592(I13462,g2380,g2384);
  nand NAND_17593(I13463,g2380,I13462);
  nand NAND_17594(I13464,g2384,I13462);
  nand NAND_17595(g9912,I13463,I13464);
  nand NAND_17596(g9954,g6128,g6120);
  nand NAND_17597(I13497,g255,g232);
  nand NAND_17598(I13498,g255,I13497);
  nand NAND_17599(I13499,g232,I13497);
  nand NAND_17600(g9966,I13498,I13499);
  nand NAND_17601(I13509,g2089,g2093);
  nand NAND_17602(I13510,g2089,I13509);
  nand NAND_17603(I13511,g2093,I13509);
  nand NAND_17604(g9972,I13510,I13511);
  nand NAND_17605(I13518,g2514,g2518);
  nand NAND_17606(I13519,g2514,I13518);
  nand NAND_17607(I13520,g2518,I13518);
  nand NAND_17608(g9975,I13519,I13520);
  nand NAND_17609(g10022,g6474,g6466);
  nand NAND_17610(I13564,g2648,g2652);
  nand NAND_17611(I13565,g2648,I13564);
  nand NAND_17612(I13566,g2652,I13564);
  nand NAND_17613(g10041,I13565,I13566);
  nand NAND_17614(g10124,g5276,g5320,g5290,g5313);
  nand NAND_17615(g10160,g5623,g5666,g5637,g5659);
  nand NAND_17616(g10185,g5969,g6012,g5983,g6005);
  nand NAND_17617(g10207,g6315,g6358,g6329,g6351);
  nand NAND_17618(g10224,g6661,g6704,g6675,g6697);
  nand NAND_17619(I13729,g4534,g4537);
  nand NAND_17620(I13730,g4534,I13729);
  nand NAND_17621(I13731,g4537,I13729);
  nand NAND_17622(g10307,I13730,I13731);
  nand NAND_17623(I13749,g4608,g4584);
  nand NAND_17624(I13750,g4608,I13749);
  nand NAND_17625(I13751,g4584,I13749);
  nand NAND_17626(g10336,I13750,I13751);
  nand NAND_17627(I13850,g862,g7397);
  nand NAND_17628(I13851,g862,I13850);
  nand NAND_17629(I13852,g7397,I13850);
  nand NAND_17630(g10472,I13851,I13852);
  nand NAND_17631(g10511,g4628,g7202,g4621);
  nand NAND_17632(g10515,g10337,g5022);
  nand NAND_17633(g10520,g7195,g7115);
  nand NAND_17634(g10529,g1592,g7308);
  nand NAND_17635(g10537,g7138,g5366);
  nand NAND_17636(g10550,g7268,g7308);
  nand NAND_17637(g10551,g1728,g7356);
  nand NAND_17638(g10552,g2153,g7374);
  nand NAND_17639(g10556,g7971,g8133);
  nand NAND_17640(g10561,g7157,g5712);
  nand NAND_17641(g10566,g7315,g7356);
  nand NAND_17642(g10567,g1862,g7405);
  nand NAND_17643(g10568,g7328,g7374);
  nand NAND_17644(g10569,g2287,g7418);
  nand NAND_17645(g10573,g7992,g8179);
  nand NAND_17646(g10578,g7174,g6058);
  nand NAND_17647(g10583,g7475,g862);
  nand NAND_17648(g10584,g7362,g7405);
  nand NAND_17649(g10585,g1996,g7451);
  nand NAND_17650(g10586,g7380,g7418);
  nand NAND_17651(g10587,g2421,g7456);
  nand NAND_17652(g10598,g7191,g6404);
  nand NAND_17653(g10601,g896,g7397);
  nand NAND_17654(g10602,g7411,g7451);
  nand NAND_17655(g10603,g10077,g9751);
  nand NAND_17656(g10604,g7424,g7456);
  nand NAND_17657(g10605,g2555,g7490);
  nand NAND_17658(g10609,g10111,g9826);
  nand NAND_17659(g10610,g7462,g7490);
  nand NAND_17660(g10611,g10115,g9831);
  nand NAND_17661(g10614,g9024,g8977,g8928);
  nand NAND_17662(g10617,g10151,g9909);
  nand NAND_17663(g10618,g10153,g9913);
  nand NAND_17664(g10622,g10178,g9973);
  nand NAND_17665(g10623,g10181,g9976);
  nand NAND_17666(g10653,g10204,g10042);
  nand NAND_17667(g10726,g7304,g7661,g979,g1061);
  nand NAND_17668(g10737,g6961,g9848);
  nand NAND_17669(g10738,g6961,g10308);
  nand NAND_17670(g10754,g7936,g7913,g8411);
  nand NAND_17671(g10755,g7352,g7675,g1322,g1404);
  nand NAND_17672(g10759,g7537,g324);
  nand NAND_17673(g10775,g7960,g7943,g8470);
  nand NAND_17674(g10796,g7537,g7523);
  nand NAND_17675(g10820,g9985,g9920,g9843);
  nand NAND_17676(g10905,g1116,g7304);
  nand NAND_17677(g10909,g7304,g1116);
  nand NAND_17678(g10916,g1146,g7854);
  nand NAND_17679(g10928,g8181,g8137,g417);
  nand NAND_17680(g10929,g1099,g7854);
  nand NAND_17681(g10935,g1459,g7352);
  nand NAND_17682(g10939,g7352,g1459);
  nand NAND_17683(g10946,g1489,g7876);
  nand NAND_17684(g10951,g7845,g7868);
  nand NAND_17685(g10961,g1442,g7876);
  nand NAND_17686(g10971,g7867,g7886);
  nand NAND_17687(g11002,g7475,g862);
  nand NAND_17688(g11020,g9187,g9040);
  nand NAND_17689(g11117,g8087,g8186,g8239);
  nand NAND_17690(I14169,g8389,g3119);
  nand NAND_17691(I14170,g8389,I14169);
  nand NAND_17692(I14171,g3119,I14169);
  nand NAND_17693(g11118,I14170,I14171);
  nand NAND_17694(g11130,g1221,g7918);
  nand NAND_17695(g11134,g8138,g8240,g8301);
  nand NAND_17696(I14185,g8442,g3470);
  nand NAND_17697(I14186,g8442,I14185);
  nand NAND_17698(I14187,g3470,I14185);
  nand NAND_17699(g11135,I14186,I14187);
  nand NAND_17700(g11149,g1564,g7948);
  nand NAND_17701(I14204,g8508,g3821);
  nand NAND_17702(I14205,g8508,I14204);
  nand NAND_17703(I14206,g3821,I14204);
  nand NAND_17704(g11153,I14205,I14206);
  nand NAND_17705(I14211,g9252,g9295);
  nand NAND_17706(I14212,g9252,I14211);
  nand NAND_17707(I14213,g9295,I14211);
  nand NAND_17708(g11154,I14212,I14213);
  nand NAND_17709(g11155,g4776,g7892,g9030);
  nand NAND_17710(I14228,g979,g8055);
  nand NAND_17711(I14229,g979,I14228);
  nand NAND_17712(I14230,g8055,I14228);
  nand NAND_17713(g11169,I14229,I14230);
  nand NAND_17714(g11172,g8478,g3096);
  nand NAND_17715(g11173,g4966,g7898,g9064);
  nand NAND_17716(I14247,g1322,g8091);
  nand NAND_17717(I14248,g1322,I14247);
  nand NAND_17718(I14249,g8091,I14247);
  nand NAND_17719(g11189,I14248,I14249);
  nand NAND_17720(g11190,g8539,g3447);
  nand NAND_17721(I14257,g8154,g3133);
  nand NAND_17722(I14258,g8154,I14257);
  nand NAND_17723(I14259,g3133,I14257);
  nand NAND_17724(g11193,I14258,I14259);
  nand NAND_17725(g11200,g8592,g3798);
  nand NAND_17726(I14275,g8218,g3484);
  nand NAND_17727(I14276,g8218,I14275);
  nand NAND_17728(I14277,g3484,I14275);
  nand NAND_17729(g11206,I14276,I14277);
  nand NAND_17730(I14289,g8282,g3835);
  nand NAND_17731(I14290,g8282,I14289);
  nand NAND_17732(I14291,g3835,I14289);
  nand NAND_17733(g11224,I14290,I14291);
  nand NAND_17734(g11245,g7636,g7733,g7697);
  nand NAND_17735(g11251,g8438,g3092);
  nand NAND_17736(g11279,g8504,g3443);
  nand NAND_17737(I14330,g225,g9966);
  nand NAND_17738(I14331,g225,I14330);
  nand NAND_17739(I14332,g9966,I14330);
  nand NAND_17740(g11292,I14331,I14332);
  nand NAND_17741(g11302,g9496,g3281);
  nand NAND_17742(g11312,g8565,g3794);
  nand NAND_17743(g11320,g4633,g4621,g7202);
  nand NAND_17744(I14350,g8890,g8848);
  nand NAND_17745(I14351,g8890,I14350);
  nand NAND_17746(I14352,g8848,I14350);
  nand NAND_17747(g11323,I14351,I14352);
  nand NAND_17748(g11326,g8993,g376,g365,g370);
  nand NAND_17749(g11330,g9483,g1193);
  nand NAND_17750(I14368,g8481,g3303);
  nand NAND_17751(I14369,g8481,I14368);
  nand NAND_17752(I14370,g3303,I14368);
  nand NAND_17753(g11350,I14369,I14370);
  nand NAND_17754(g11355,g9551,g3310);
  nand NAND_17755(g11356,g9552,g3632);
  nand NAND_17756(g11374,g9536,g1536);
  nand NAND_17757(g11381,g9660,g3274);
  nand NAND_17758(g11382,g8644,g6895,g8663);
  nand NAND_17759(I14398,g8542,g3654);
  nand NAND_17760(I14399,g8542,I14398);
  nand NAND_17761(I14400,g3654,I14398);
  nand NAND_17762(g11389,I14399,I14400);
  nand NAND_17763(g11394,g9600,g3661);
  nand NAND_17764(g11395,g9601,g3983);
  nand NAND_17765(g11396,g8713,g4688);
  nand NAND_17766(g11405,g2741,g2735,g6856,g2748);
  nand NAND_17767(g11409,g9842,g3298);
  nand NAND_17768(g11410,g6875,g6895,g8696);
  nand NAND_17769(g11411,g9713,g3625);
  nand NAND_17770(g11412,g8666,g6918,g8697);
  nand NAND_17771(I14427,g8595,g4005);
  nand NAND_17772(I14428,g8595,I14427);
  nand NAND_17773(I14429,g4005,I14427);
  nand NAND_17774(g11419,I14428,I14429);
  nand NAND_17775(g11424,g9662,g4012);
  nand NAND_17776(g11426,g8742,g4878);
  nand NAND_17777(g11432,g10295,g8864);
  nand NAND_17778(g11441,g9599,g3267);
  nand NAND_17779(g11442,g8644,g3288,g3343);
  nand NAND_17780(g11443,g9916,g3649);
  nand NAND_17781(g11444,g6905,g6918,g8733);
  nand NAND_17782(g11445,g9771,g3976);
  nand NAND_17783(g11446,g8700,g6941,g8734);
  nand NAND_17784(g11479,g6875,g3288,g3347);
  nand NAND_17785(g11480,g10323,g8906);
  nand NAND_17786(g11489,g9661,g3618);
  nand NAND_17787(g11490,g8666,g3639,g3694);
  nand NAND_17788(g11491,g9982,g4000);
  nand NAND_17789(g11492,g6928,g6941,g8756);
  nand NAND_17790(I14480,g10074,g655);
  nand NAND_17791(I14481,g10074,I14480);
  nand NAND_17792(I14482,g655,I14480);
  nand NAND_17793(g11511,I14481,I14482);
  nand NAND_17794(g11533,g6905,g3639,g3698);
  nand NAND_17795(g11534,g7121,g8958);
  nand NAND_17796(g11543,g9714,g3969);
  nand NAND_17797(g11544,g8700,g3990,g4045);
  nand NAND_17798(I14497,g9020,g8737);
  nand NAND_17799(I14498,g9020,I14497);
  nand NAND_17800(I14499,g8737,I14497);
  nand NAND_17801(g11545,I14498,I14499);
  nand NAND_17802(I14508,g370,g8721);
  nand NAND_17803(I14509,g370,I14508);
  nand NAND_17804(I14510,g8721,I14508);
  nand NAND_17805(g11559,I14509,I14510);
  nand NAND_17806(I14516,g10147,g661);
  nand NAND_17807(I14517,g10147,I14516);
  nand NAND_17808(I14518,g661,I14516);
  nand NAND_17809(g11561,I14517,I14518);
  nand NAND_17810(g11590,g6928,g3990,g4049);
  nand NAND_17811(I14530,g8840,g8873);
  nand NAND_17812(I14531,g8840,I14530);
  nand NAND_17813(I14532,g8873,I14530);
  nand NAND_17814(g11591,I14531,I14532);
  nand NAND_17815(g11639,g8933,g4722);
  nand NAND_17816(g11674,g8676,g4674);
  nand NAND_17817(g11675,g8984,g4912);
  nand NAND_17818(g11676,g358,g8944,g376,g385);
  nand NAND_17819(g11679,g8836,g802);
  nand NAND_17820(g11707,g8718,g4864);
  nand NAND_17821(g11708,g10147,g10110);
  nand NAND_17822(I14609,g8993,g8678);
  nand NAND_17823(I14610,g8993,I14609);
  nand NAND_17824(I14611,g8678,I14609);
  nand NAND_17825(g11761,I14610,I14611);
  nand NAND_17826(g11858,g9014,g3010);
  nand NAND_17827(g11881,g9060,g3361);
  nand NAND_17828(g11892,g7777,g9086);
  nand NAND_17829(g11903,g9099,g3712);
  nand NAND_17830(I14712,g9671,g5128);
  nand NAND_17831(I14713,g9671,I14712);
  nand NAND_17832(I14714,g5128,I14712);
  nand NAND_17833(g11906,I14713,I14714);
  nand NAND_17834(g11914,g8187,g1648);
  nand NAND_17835(I14733,g9732,g5475);
  nand NAND_17836(I14734,g9732,I14733);
  nand NAND_17837(I14735,g5475,I14733);
  nand NAND_17838(g11923,I14734,I14735);
  nand NAND_17839(g11933,g837,g9334,g7197);
  nand NAND_17840(g11934,g8139,g8187);
  nand NAND_17841(g11936,g8241,g1783);
  nand NAND_17842(g11938,g8259,g2208);
  nand NAND_17843(I14764,g9808,g5821);
  nand NAND_17844(I14765,g9808,I14764);
  nand NAND_17845(I14766,g5821,I14764);
  nand NAND_17846(g11944,I14765,I14766);
  nand NAND_17847(g11951,g9166,g847,g703);
  nand NAND_17848(g11952,g1624,g8187);
  nand NAND_17849(g11953,g8195,g8241);
  nand NAND_17850(g11955,g8302,g1917);
  nand NAND_17851(g11957,g8205,g8259);
  nand NAND_17852(g11959,g8316,g2342);
  nand NAND_17853(g11961,g9777,g5105);
  nand NAND_17854(I14788,g9891,g6167);
  nand NAND_17855(I14789,g9891,I14788);
  nand NAND_17856(I14790,g6167,I14788);
  nand NAND_17857(g11962,I14789,I14790);
  nand NAND_17858(g11968,g837,g9334,g9086);
  nand NAND_17859(g11969,g7252,g1636);
  nand NAND_17860(g11970,g1760,g8241);
  nand NAND_17861(g11971,g8249,g8302);
  nand NAND_17862(g11973,g8365,g2051);
  nand NAND_17863(g11974,g2185,g8259);
  nand NAND_17864(g11975,g8267,g8316);
  nand NAND_17865(g11977,g8373,g2476);
  nand NAND_17866(g11979,g9861,g5452);
  nand NAND_17867(I14816,g9962,g6513);
  nand NAND_17868(I14817,g9962,I14816);
  nand NAND_17869(I14818,g6513,I14816);
  nand NAND_17870(g11980,I14817,I14818);
  nand NAND_17871(g11990,g9166,g703);
  nand NAND_17872(g11992,g7275,g1772);
  nand NAND_17873(g11993,g1894,g8302);
  nand NAND_17874(g11994,g8310,g8365);
  nand NAND_17875(g11996,g7280,g2197);
  nand NAND_17876(g11997,g2319,g8316);
  nand NAND_17877(g11998,g8324,g8373);
  nand NAND_17878(g12000,g8418,g2610);
  nand NAND_17879(I14853,g9433,g5142);
  nand NAND_17880(I14854,g9433,I14853);
  nand NAND_17881(I14855,g5142,I14853);
  nand NAND_17882(g12001,I14854,I14855);
  nand NAND_17883(g12008,g9932,g5798);
  nand NAND_17884(g12014,g7197,g703);
  nand NAND_17885(g12016,g1648,g8093);
  nand NAND_17886(g12019,g7322,g1906);
  nand NAND_17887(g12020,g2028,g8365);
  nand NAND_17888(g12022,g7335,g2331);
  nand NAND_17889(g12023,g2453,g8373);
  nand NAND_17890(g12024,g8381,g8418);
  nand NAND_17891(I14883,g9500,g5489);
  nand NAND_17892(I14884,g9500,I14883);
  nand NAND_17893(I14885,g5489,I14883);
  nand NAND_17894(g12028,I14884,I14885);
  nand NAND_17895(g12035,g10000,g6144);
  nand NAND_17896(g12042,g9086,g703);
  nand NAND_17897(g12044,g1657,g8139);
  nand NAND_17898(g12045,g1783,g8146);
  nand NAND_17899(g12048,g7369,g2040);
  nand NAND_17900(g12049,g2208,g8150);
  nand NAND_17901(g12052,g7387,g2465);
  nand NAND_17902(g12053,g2587,g8418);
  nand NAND_17903(I14923,g9558,g5835);
  nand NAND_17904(I14924,g9558,I14923);
  nand NAND_17905(I14925,g5835,I14923);
  nand NAND_17906(g12066,I14924,I14925);
  nand NAND_17907(g12073,g10058,g6490);
  nand NAND_17908(g12078,g8187,g8093);
  nand NAND_17909(g12079,g1792,g8195);
  nand NAND_17910(g12080,g1917,g8201);
  nand NAND_17911(g12083,g2217,g8205);
  nand NAND_17912(g12084,g2342,g8211);
  nand NAND_17913(g12087,g7431,g2599);
  nand NAND_17914(I14955,g9620,g6181);
  nand NAND_17915(I14956,g9620,I14955);
  nand NAND_17916(I14957,g6181,I14955);
  nand NAND_17917(g12100,I14956,I14957);
  nand NAND_17918(g12111,g847,g9166);
  nand NAND_17919(g12112,g8139,g1624);
  nand NAND_17920(g12114,g8241,g8146);
  nand NAND_17921(g12115,g1926,g8249);
  nand NAND_17922(g12116,g2051,g8255);
  nand NAND_17923(g12118,g8259,g8150);
  nand NAND_17924(g12119,g2351,g8267);
  nand NAND_17925(g12120,g2476,g8273);
  nand NAND_17926(g12124,g8741,g4674);
  nand NAND_17927(g12125,g9728,g5101);
  nand NAND_17928(I14991,g9685,g6527);
  nand NAND_17929(I14992,g9685,I14991);
  nand NAND_17930(I14993,g6527,I14991);
  nand NAND_17931(g12136,I14992,I14993);
  nand NAND_17932(I15002,g9691,g1700);
  nand NAND_17933(I15003,g9691,I15002);
  nand NAND_17934(I15004,g1700,I15002);
  nand NAND_17935(g12144,I15003,I15004);
  nand NAND_17936(g12145,g8195,g1760);
  nand NAND_17937(g12147,g8302,g8201);
  nand NAND_17938(g12148,g2060,g8310);
  nand NAND_17939(g12149,g8205,g2185);
  nand NAND_17940(g12151,g8316,g8211);
  nand NAND_17941(g12152,g2485,g8324);
  nand NAND_17942(g12153,g2610,g8330);
  nand NAND_17943(g12155,g7753,g7717);
  nand NAND_17944(g12159,g8765,g4864);
  nand NAND_17945(g12169,g9804,g5448);
  nand NAND_17946(g12185,g9905,g799);
  nand NAND_17947(I15041,g9752,g1834);
  nand NAND_17948(I15042,g9752,I15041);
  nand NAND_17949(I15043,g1834,I15041);
  nand NAND_17950(g12187,I15042,I15043);
  nand NAND_17951(g12188,g8249,g1894);
  nand NAND_17952(g12190,g8365,g8255);
  nand NAND_17953(I15051,g9759,g2259);
  nand NAND_17954(I15052,g9759,I15051);
  nand NAND_17955(I15053,g2259,I15051);
  nand NAND_17956(g12191,I15052,I15053);
  nand NAND_17957(g12192,g8267,g2319);
  nand NAND_17958(g12194,g8373,g8273);
  nand NAND_17959(g12195,g2619,g8381);
  nand NAND_17960(g12196,g8764,g4688);
  nand NAND_17961(g12197,g7296,g5290);
  nand NAND_17962(g12207,g9887,g5794);
  nand NAND_17963(I15078,g9827,g1968);
  nand NAND_17964(I15079,g9827,I15078);
  nand NAND_17965(I15080,g1968,I15078);
  nand NAND_17966(g12221,I15079,I15080);
  nand NAND_17967(g12222,g8310,g2028);
  nand NAND_17968(I15087,g9832,g2393);
  nand NAND_17969(I15088,g9832,I15087);
  nand NAND_17970(I15089,g2393,I15087);
  nand NAND_17971(g12224,I15088,I15089);
  nand NAND_17972(g12225,g8324,g2453);
  nand NAND_17973(g12227,g8418,g8330);
  nand NAND_17974(g12232,g8804,g4878);
  nand NAND_17975(I15105,g9780,g5313);
  nand NAND_17976(I15106,g9780,I15105);
  nand NAND_17977(I15107,g5313,I15105);
  nand NAND_17978(g12239,I15106,I15107);
  nand NAND_17979(g12244,g7343,g5320);
  nand NAND_17980(g12245,g7344,g5637);
  nand NAND_17981(g12255,g9958,g6140);
  nand NAND_17982(I15121,g9910,g2102);
  nand NAND_17983(I15122,g9910,I15121);
  nand NAND_17984(I15123,g2102,I15121);
  nand NAND_17985(g12285,I15122,I15123);
  nand NAND_17986(I15128,g9914,g2527);
  nand NAND_17987(I15129,g9914,I15128);
  nand NAND_17988(I15130,g2527,I15128);
  nand NAND_17989(g12286,I15129,I15130);
  nand NAND_17990(g12287,g8381,g2587);
  nand NAND_17991(g12289,g9978,g9766,g9708);
  nand NAND_17992(g12292,g4698,g8933);
  nand NAND_17993(g12293,g7436,g5283);
  nand NAND_17994(g12294,g10044,g7018,g10090);
  nand NAND_17995(I15147,g9864,g5659);
  nand NAND_17996(I15148,g9864,I15147);
  nand NAND_17997(I15149,g5659,I15147);
  nand NAND_17998(g12301,I15148,I15149);
  nand NAND_17999(g12306,g7394,g5666);
  nand NAND_18000(g12307,g7395,g5983);
  nand NAND_18001(g12317,g10026,g6486);
  nand NAND_18002(g12323,g9480,g640);
  nand NAND_18003(I15166,g9904,g9823);
  nand NAND_18004(I15167,g9904,I15166);
  nand NAND_18005(I15168,g9823,I15166);
  nand NAND_18006(g12332,I15167,I15168);
  nand NAND_18007(I15174,g9977,g2661);
  nand NAND_18008(I15175,g9977,I15174);
  nand NAND_18009(I15176,g2661,I15174);
  nand NAND_18010(g12336,I15175,I15176);
  nand NAND_18011(g12340,g4888,g8984);
  nand NAND_18012(g12341,g7512,g5308);
  nand NAND_18013(g12342,g7004,g7018,g10129);
  nand NAND_18014(g12343,g7470,g5630);
  nand NAND_18015(g12344,g10093,g7041,g10130);
  nand NAND_18016(I15193,g9935,g6005);
  nand NAND_18017(I15194,g9935,I15193);
  nand NAND_18018(I15195,g6005,I15193);
  nand NAND_18019(g12351,I15194,I15195);
  nand NAND_18020(g12356,g7438,g6012);
  nand NAND_18021(g12357,g7439,g6329);
  nand NAND_18022(g12369,g9049,g637);
  nand NAND_18023(I15212,g10035,g1714);
  nand NAND_18024(I15213,g10035,I15212);
  nand NAND_18025(I15214,g1714,I15212);
  nand NAND_18026(g12370,I15213,I15214);
  nand NAND_18027(g12402,g7704,g10266);
  nand NAND_18028(g12411,g7393,g5276);
  nand NAND_18029(g12412,g10044,g5297,g5348);
  nand NAND_18030(g12413,g7521,g5654);
  nand NAND_18031(g12414,g7028,g7041,g10165);
  nand NAND_18032(g12415,g7496,g5976);
  nand NAND_18033(g12416,g10133,g7064,g10166);
  nand NAND_18034(I15241,g10003,g6351);
  nand NAND_18035(I15242,g10003,I15241);
  nand NAND_18036(I15243,g6351,I15241);
  nand NAND_18037(g12423,I15242,I15243);
  nand NAND_18038(g12428,g7472,g6358);
  nand NAND_18039(g12429,g7473,g6675);
  nand NAND_18040(I15253,g10078,g1848);
  nand NAND_18041(I15254,g10078,I15253);
  nand NAND_18042(I15255,g1848,I15253);
  nand NAND_18043(g12431,I15254,I15255);
  nand NAND_18044(I15262,g10081,g2273);
  nand NAND_18045(I15263,g10081,I15262);
  nand NAND_18046(I15264,g2273,I15262);
  nand NAND_18047(g12436,I15263,I15264);
  nand NAND_18048(g12449,g7004,g5297,g5352);
  nand NAND_18049(g12450,g7738,g10281);
  nand NAND_18050(g12459,g7437,g5623);
  nand NAND_18051(g12460,g10093,g5644,g5694);
  nand NAND_18052(g12461,g7536,g6000);
  nand NAND_18053(g12462,g7051,g7064,g10190);
  nand NAND_18054(g12463,g7513,g6322);
  nand NAND_18055(g12464,g10169,g7087,g10191);
  nand NAND_18056(I15287,g10061,g6697);
  nand NAND_18057(I15288,g10061,I15287);
  nand NAND_18058(I15289,g6697,I15287);
  nand NAND_18059(g12471,I15288,I15289);
  nand NAND_18060(g12476,g7498,g6704);
  nand NAND_18061(I15298,g10112,g1982);
  nand NAND_18062(I15299,g10112,I15298);
  nand NAND_18063(I15300,g1982,I15298);
  nand NAND_18064(g12478,I15299,I15300);
  nand NAND_18065(I15306,g10116,g2407);
  nand NAND_18066(I15307,g10116,I15306);
  nand NAND_18067(I15308,g2407,I15306);
  nand NAND_18068(g12482,I15307,I15308);
  nand NAND_18069(g12491,g7285,g4462,g6961);
  nand NAND_18070(g12511,g7028,g5644,g5698);
  nand NAND_18071(g12512,g7766,g10312);
  nand NAND_18072(g12521,g7471,g5969);
  nand NAND_18073(g12522,g10133,g5990,g6040);
  nand NAND_18074(g12523,g7563,g6346);
  nand NAND_18075(g12524,g7074,g7087,g10212);
  nand NAND_18076(g12525,g7522,g6668);
  nand NAND_18077(g12526,g10194,g7110,g10213);
  nand NAND_18078(I15333,g10152,g2116);
  nand NAND_18079(I15334,g10152,I15333);
  nand NAND_18080(I15335,g2116,I15333);
  nand NAND_18081(g12538,I15334,I15335);
  nand NAND_18082(I15340,g10154,g2541);
  nand NAND_18083(I15341,g10154,I15340);
  nand NAND_18084(I15342,g2541,I15340);
  nand NAND_18085(g12539,I15341,I15342);
  nand NAND_18086(g12577,g7051,g5990,g6044);
  nand NAND_18087(g12578,g7791,g10341);
  nand NAND_18088(g12587,g7497,g6315);
  nand NAND_18089(g12588,g10169,g6336,g6386);
  nand NAND_18090(g12589,g7591,g6692);
  nand NAND_18091(g12590,g7097,g7110,g10229);
  nand NAND_18092(I15363,g10182,g2675);
  nand NAND_18093(I15364,g10182,I15363);
  nand NAND_18094(I15365,g2675,I15363);
  nand NAND_18095(g12592,I15364,I15365);
  nand NAND_18096(g12628,g7074,g6336,g6390);
  nand NAND_18097(g12629,g7812,g7142);
  nand NAND_18098(g12638,g7514,g6661);
  nand NAND_18099(g12639,g10194,g6682,g6732);
  nand NAND_18100(g12644,g10233,g4531);
  nand NAND_18101(g12686,g7097,g6682,g6736);
  nand NAND_18102(g12767,g4467,g6961);
  nand NAND_18103(g12796,g4467,g6961);
  nand NAND_18104(g12797,g10275,g7655,g7643,g7627);
  nand NAND_18105(g12819,g9848,g6961);
  nand NAND_18106(g12822,g6978,g7236,g7224,g7163);
  nand NAND_18107(g12910,g11002,g10601);
  nand NAND_18108(g12915,g12806,g12632);
  nand NAND_18109(g12933,g7150,g10515);
  nand NAND_18110(g12941,g7167,g10537);
  nand NAND_18111(g12947,g7184,g10561);
  nand NAND_18112(g12969,g4388,g7178,g10476);
  nand NAND_18113(g12971,g9024,g8977,g10664);
  nand NAND_18114(g12972,g7209,g10578);
  nand NAND_18115(g12999,g4392,g10476,g4401);
  nand NAND_18116(g13000,g7228,g10598);
  nand NAND_18117(g13040,g5196,g12002,g5308,g9780);
  nand NAND_18118(g13043,g10521,g969);
  nand NAND_18119(g13050,g5543,g12029,g5654,g9864);
  nand NAND_18120(g13057,g969,g11294);
  nand NAND_18121(g13058,g10544,g1312);
  nand NAND_18122(g13066,g4430,g7178,g10590);
  nand NAND_18123(g13067,g5240,g12059,g5331,g9780);
  nand NAND_18124(g13069,g5889,g12067,g6000,g9935);
  nand NAND_18125(g13079,g1312,g11336);
  nand NAND_18126(g13083,g4392,g10590,g4434);
  nand NAND_18127(g13084,g5587,g12093,g5677,g9864);
  nand NAND_18128(g13086,g6235,g12101,g6346,g10003);
  nand NAND_18129(g13092,g1061,g10761);
  nand NAND_18130(g13093,g10649,g7661,g979,g1061);
  nand NAND_18131(g13097,g5204,g12002,g5339,g9780);
  nand NAND_18132(g13098,g5933,g12129,g6023,g9935);
  nand NAND_18133(g13100,g6581,g12137,g6692,g10061);
  nand NAND_18134(g13102,g7523,g10759);
  nand NAND_18135(g13104,g1404,g10794);
  nand NAND_18136(g13105,g10671,g7675,g1322,g1404);
  nand NAND_18137(g13108,g5551,g12029,g5685,g9864);
  nand NAND_18138(g13109,g6279,g12173,g6369,g10003);
  nand NAND_18139(g13115,g1008,g11786,g11294);
  nand NAND_18140(g13118,g5897,g12067,g6031,g9935);
  nand NAND_18141(g13119,g6625,g12211,g6715,g10061);
  nand NAND_18142(g13121,g11117,g8411);
  nand NAND_18143(g13124,g10666,g7661,g979,g1061);
  nand NAND_18144(g13130,g1351,g11815,g11336);
  nand NAND_18145(g13131,g6243,g12101,g6377,g10003);
  nand NAND_18146(g13134,g11134,g8470);
  nand NAND_18147(g13137,g10699,g7675,g1322,g1404);
  nand NAND_18148(g13139,g6589,g12137,g6723,g10061);
  nand NAND_18149(g13143,g10695,g7661,g979,g1061);
  nand NAND_18150(g13176,g10715,g7675,g1322,g1404);
  nand NAND_18151(g13210,g7479,g10521);
  nand NAND_18152(g13217,g4082,g10808);
  nand NAND_18153(g13240,g1046,g10521);
  nand NAND_18154(g13241,g7503,g10544);
  nand NAND_18155(g13248,g9985,g12399,g9843);
  nand NAND_18156(g13256,g11846,g11294,g11812);
  nand NAND_18157(g13257,g1389,g10544);
  nand NAND_18158(g13260,g1116,g10666);
  nand NAND_18159(g13264,g11869,g11336,g11849);
  nand NAND_18160(g13266,g12440,g9920,g9843);
  nand NAND_18161(g13273,g1459,g10699);
  nand NAND_18162(g13281,g10916,g1099);
  nand NAND_18163(g13283,g12440,g12399,g9843);
  nand NAND_18164(g13284,g10695,g1157);
  nand NAND_18165(g13288,g10946,g1442);
  nand NAND_18166(g13291,g10715,g1500);
  nand NAND_18167(g13307,g1116,g10695);
  nand NAND_18168(g13315,g1459,g10715);
  nand NAND_18169(g13330,g4664,g11006);
  nand NAND_18170(g13346,g4854,g11012);
  nand NAND_18171(g13432,g4793,g10831);
  nand NAND_18172(g13459,g7479,g11294,g11846);
  nand NAND_18173(g13462,g12449,g12412,g12342,g12294);
  nand NAND_18174(g13464,g10831,g4793,g4776);
  nand NAND_18175(g13469,g4983,g10862);
  nand NAND_18176(g13475,g1008,g11294,g11786);
  nand NAND_18177(g13476,g7503,g11336,g11869);
  nand NAND_18178(g13478,g12511,g12460,g12414,g12344);
  nand NAND_18179(g13479,g12686,g12639,g12590,g12526);
  nand NAND_18180(g13486,g10862,g4983,g4966);
  nand NAND_18181(g13495,g1008,g11786,g7972);
  nand NAND_18182(g13496,g1351,g11336,g11815);
  nand NAND_18183(g13498,g12577,g12522,g12462,g12416);
  nand NAND_18184(g13499,g11479,g11442,g11410,g11382);
  nand NAND_18185(g13511,g182,g174,g203,g12812);
  nand NAND_18186(g13513,g1351,g11815,g8002);
  nand NAND_18187(g13515,g12628,g12588,g12524,g12464);
  nand NAND_18188(g13516,g11533,g11490,g11444,g11412);
  nand NAND_18189(g13527,g182,g168,g203,g12812);
  nand NAND_18190(g13528,g11294,g7549,g1008);
  nand NAND_18191(g13529,g11590,g11544,g11492,g11446);
  nand NAND_18192(g13544,g7972,g10521,g7549,g1008);
  nand NAND_18193(g13551,g11812,g7479,g7903,g10521);
  nand NAND_18194(g13554,g11336,g7582,g1351);
  nand NAND_18195(g13573,g8002,g10544,g7582,g1351);
  nand NAND_18196(g13580,g11849,g7503,g7922,g10544);
  nand NAND_18197(g13600,g3021,g11039);
  nand NAND_18198(g13627,g11172,g8388);
  nand NAND_18199(g13628,g3372,g11107);
  nand NAND_18200(g13634,g11797,g11261);
  nand NAND_18201(g13666,g11190,g8441);
  nand NAND_18202(g13667,g3723,g11119);
  nand NAND_18203(g13672,g8933,g11261);
  nand NAND_18204(g13676,g11834,g11283);
  nand NAND_18205(g13708,g11200,g8507);
  nand NAND_18206(g13709,g11755,g11261);
  nand NAND_18207(g13712,g8984,g11283);
  nand NAND_18208(g13727,g174,g203,g168,g12812);
  nand NAND_18209(g13739,g11773,g11261);
  nand NAND_18210(g13742,g11780,g11283);
  nand NAND_18211(g13756,g203,g12812);
  nand NAND_18212(g13764,g11252,g3072);
  nand NAND_18213(g13779,g11804,g11283);
  nand NAND_18214(g13795,g11216,g401);
  nand NAND_18215(g13797,g8102,g11273);
  nand NAND_18216(g13798,g11280,g3423);
  nand NAND_18217(g13821,g11251,g8340);
  nand NAND_18218(g13822,g8160,g11306);
  nand NAND_18219(g13823,g11313,g3774);
  nand NAND_18220(g13834,g4754,g11773);
  nand NAND_18221(g13846,g1116,g10649);
  nand NAND_18222(g13850,g11279,g8396);
  nand NAND_18223(g13851,g8224,g11360);
  nand NAND_18224(g13854,g4765,g11797);
  nand NAND_18225(g13855,g4944,g11804);
  nand NAND_18226(g13861,g1459,g10671);
  nand NAND_18227(g13866,g3239,g11194,g3321,g11519);
  nand NAND_18228(g13867,g11312,g8449);
  nand NAND_18229(g13870,g11773,g4732);
  nand NAND_18230(g13871,g4955,g11834);
  nand NAND_18231(g13873,g11566,g11729);
  nand NAND_18232(g13882,g3590,g11207,g3672,g11576);
  nand NAND_18233(g13884,g11797,g4727);
  nand NAND_18234(g13886,g11804,g4922);
  nand NAND_18235(g13889,g11566,g11435);
  nand NAND_18236(g13892,g11653,g11473);
  nand NAND_18237(g13896,g3227,g11194,g3281,g11350);
  nand NAND_18238(g13897,g3211,g11217,g3329,g11519);
  nand NAND_18239(g13898,g11621,g11747);
  nand NAND_18240(g13907,g3941,g11225,g4023,g11631);
  nand NAND_18241(g13909,g11396,g8847,g11674,g8803);
  nand NAND_18242(g13911,g11834,g4917);
  nand NAND_18243(g13915,g11566,g11473);
  nand NAND_18244(g13918,g3259,g11217,g3267,g11350);
  nand NAND_18245(g13920,g11621,g11483);
  nand NAND_18246(g13923,g11692,g11527);
  nand NAND_18247(g13927,g3578,g11207,g3632,g11389);
  nand NAND_18248(g13928,g3562,g11238,g3680,g11576);
  nand NAND_18249(g13929,g11669,g11763);
  nand NAND_18250(g13940,g11426,g8889,g11707,g8829);
  nand NAND_18251(g13945,g691,g11740);
  nand NAND_18252(g13948,g11610,g8864);
  nand NAND_18253(g13951,g10295,g11729);
  nand NAND_18254(g13955,g11621,g11527);
  nand NAND_18255(g13958,g3610,g11238,g3618,g11389);
  nand NAND_18256(g13960,g11669,g11537);
  nand NAND_18257(g13963,g11715,g11584);
  nand NAND_18258(g13967,g3929,g11225,g3983,g11419);
  nand NAND_18259(g13968,g3913,g11255,g4031,g11631);
  nand NAND_18260(g13977,g11610,g11729);
  nand NAND_18261(g13980,g10295,g11435);
  nand NAND_18262(g13983,g11658,g8906);
  nand NAND_18263(g13986,g10323,g11747);
  nand NAND_18264(g13990,g11669,g11584);
  nand NAND_18265(g13993,g3961,g11255,g3969,g11419);
  nand NAND_18266(g14005,g11514,g11729);
  nand NAND_18267(g14008,g11610,g11435);
  nand NAND_18268(g14011,g10295,g11473);
  nand NAND_18269(g14014,g3199,g11217,g3298,g11519);
  nand NAND_18270(g14015,g11658,g11747);
  nand NAND_18271(g14018,g10323,g11483);
  nand NAND_18272(g14021,g11697,g8958);
  nand NAND_18273(g14024,g7121,g11763);
  nand NAND_18274(g14038,g11514,g11435);
  nand NAND_18275(g14041,g11610,g11473);
  nand NAND_18276(g14045,g11571,g11747);
  nand NAND_18277(g14048,g11658,g11483);
  nand NAND_18278(g14051,g10323,g11527);
  nand NAND_18279(g14054,g3550,g11238,g3649,g11576);
  nand NAND_18280(g14055,g11697,g11763);
  nand NAND_18281(g14058,g7121,g11537);
  nand NAND_18282(g14066,g11514,g11473);
  nand NAND_18283(g14069,g11653,g8864);
  nand NAND_18284(g14072,g11571,g11483);
  nand NAND_18285(g14075,g11658,g11527);
  nand NAND_18286(g14079,g11626,g11763);
  nand NAND_18287(g14082,g11697,g11537);
  nand NAND_18288(g14085,g7121,g11584);
  nand NAND_18289(g14088,g3901,g11255,g4000,g11631);
  nand NAND_18290(g14089,g11755,g4717);
  nand NAND_18291(g14098,g11566,g8864);
  nand NAND_18292(g14101,g11653,g11729);
  nand NAND_18293(g14104,g11514,g8864);
  nand NAND_18294(g14107,g11571,g11527);
  nand NAND_18295(g14110,g11692,g8906);
  nand NAND_18296(g14113,g11626,g11537);
  nand NAND_18297(g14116,g11697,g11584);
  nand NAND_18298(g14120,g11780,g4907);
  nand NAND_18299(g14123,g10685,g10928);
  nand NAND_18300(g14127,g11653,g11435);
  nand NAND_18301(g14130,g11621,g8906);
  nand NAND_18302(g14133,g11692,g11747);
  nand NAND_18303(g14136,g11571,g8906);
  nand NAND_18304(g14139,g11626,g11584);
  nand NAND_18305(g14142,g11715,g8958);
  nand NAND_18306(g14146,g11020,g691);
  nand NAND_18307(g14151,g11692,g11483);
  nand NAND_18308(g14154,g11669,g8958);
  nand NAND_18309(g14157,g11715,g11763);
  nand NAND_18310(g14160,g11626,g8958);
  nand NAND_18311(g14170,g11715,g11537);
  nand NAND_18312(g14177,g11741,g11721,g753);
  nand NAND_18313(g14223,g9092,g11858);
  nand NAND_18314(g14234,g9177,g11881);
  nand NAND_18315(g14254,g11968,g11933,g11951);
  nand NAND_18316(g14258,g9203,g11903);
  nand NAND_18317(g14279,g12111,g9246);
  nand NAND_18318(g14317,g5033,g11862);
  nand NAND_18319(g14333,g12042,g12014,g11990,g11892);
  nand NAND_18320(g14343,g11961,g9670);
  nand NAND_18321(g14344,g5377,g11885);
  nand NAND_18322(g14378,g11979,g9731);
  nand NAND_18323(g14379,g5723,g11907);
  nand NAND_18324(g14407,g12008,g9807);
  nand NAND_18325(g14408,g6069,g11924);
  nand NAND_18326(g14422,g3187,g11194,g3298,g8481);
  nand NAND_18327(g14433,g12035,g9890);
  nand NAND_18328(g14434,g6415,g11945);
  nand NAND_18329(g14452,g3538,g11207,g3649,g8542);
  nand NAND_18330(g14489,g12126,g5084);
  nand NAND_18331(g14505,g12073,g9961);
  nand NAND_18332(g14517,g3231,g11217,g3321,g8481);
  nand NAND_18333(g14519,g3889,g11225,g4000,g8595);
  nand NAND_18334(g14520,g9369,g12163);
  nand NAND_18335(g14521,g12170,g5428);
  nand NAND_18336(g14542,g3582,g11238,g3672,g8542);
  nand NAND_18337(g14546,g12125,g9613);
  nand NAND_18338(g14547,g9439,g12201);
  nand NAND_18339(g14548,g12208,g5774);
  nand NAND_18340(g14569,g3195,g11194,g3329,g8481);
  nand NAND_18341(g14570,g3933,g11255,g4023,g8595);
  nand NAND_18342(g14572,g12169,g9678);
  nand NAND_18343(g14573,g9506,g12249);
  nand NAND_18344(g14574,g12256,g6120);
  nand NAND_18345(g14590,g3546,g11207,g3680,g8542);
  nand NAND_18346(g14596,g12196,g9775,g12124,g9663);
  nand NAND_18347(g14598,g5248,g12002,g5331,g12497);
  nand NAND_18348(g14599,g12207,g9739);
  nand NAND_18349(g14600,g9564,g12311);
  nand NAND_18350(g14601,g12318,g6466);
  nand NAND_18351(g14625,g3897,g11225,g4031,g8595);
  nand NAND_18352(g14626,g12232,g9852,g12159,g9715);
  nand NAND_18353(g14627,g12553,g12772);
  nand NAND_18354(g14636,g5595,g12029,g5677,g12563);
  nand NAND_18355(g14637,g12255,g9815);
  nand NAND_18356(g14638,g9626,g12361);
  nand NAND_18357(g14655,g4743,g11755);
  nand NAND_18358(g14656,g12553,g12405);
  nand NAND_18359(g14659,g12646,g12443);
  nand NAND_18360(g14663,g5236,g12002,g5290,g12239);
  nand NAND_18361(g14664,g5220,g12059,g5339,g12497);
  nand NAND_18362(g14665,g12604,g12798);
  nand NAND_18363(g14674,g5941,g12067,g6023,g12614);
  nand NAND_18364(g14675,g12317,g9898);
  nand NAND_18365(I16778,g11292,g12332);
  nand NAND_18366(I16779,g11292,I16778);
  nand NAND_18367(I16780,g12332,I16778);
  nand NAND_18368(g14677,I16779,I16780);
  nand NAND_18369(g14682,g4933,g11780);
  nand NAND_18370(g14683,g12553,g12443);
  nand NAND_18371(g14686,g5268,g12059,g5276,g12239);
  nand NAND_18372(g14688,g12604,g12453);
  nand NAND_18373(g14691,g12695,g12505);
  nand NAND_18374(g14695,g5583,g12029,g5637,g12301);
  nand NAND_18375(g14696,g5567,g12093,g5685,g12563);
  nand NAND_18376(g14697,g12662,g12824);
  nand NAND_18377(g14706,g6287,g12101,g6369,g12672);
  nand NAND_18378(g14720,g12593,g10266);
  nand NAND_18379(g14723,g7704,g12772);
  nand NAND_18380(g14727,g12604,g12505);
  nand NAND_18381(g14730,g5615,g12093,g5623,g12301);
  nand NAND_18382(g14732,g12662,g12515);
  nand NAND_18383(g14735,g12739,g12571);
  nand NAND_18384(g14739,g5929,g12067,g5983,g12351);
  nand NAND_18385(g14740,g5913,g12129,g6031,g12614);
  nand NAND_18386(g14741,g12711,g10421);
  nand NAND_18387(g14750,g6633,g12137,g6715,g12721);
  nand NAND_18388(g14755,g12593,g12772);
  nand NAND_18389(g14758,g7704,g12405);
  nand NAND_18390(g14761,g12651,g10281);
  nand NAND_18391(g14764,g7738,g12798);
  nand NAND_18392(g14768,g12662,g12571);
  nand NAND_18393(g14771,g5961,g12129,g5969,g12351);
  nand NAND_18394(g14773,g12711,g12581);
  nand NAND_18395(g14776,g12780,g12622);
  nand NAND_18396(g14780,g6275,g12101,g6329,g12423);
  nand NAND_18397(g14781,g6259,g12173,g6377,g12672);
  nand NAND_18398(g14782,g12755,g10491);
  nand NAND_18399(g14794,g12492,g12772);
  nand NAND_18400(g14797,g12593,g12405);
  nand NAND_18401(g14800,g7704,g12443);
  nand NAND_18402(g14803,g5208,g12059,g5308,g12497);
  nand NAND_18403(g14804,g12651,g12798);
  nand NAND_18404(g14807,g7738,g12453);
  nand NAND_18405(g14810,g12700,g10312);
  nand NAND_18406(g14813,g7766,g12824);
  nand NAND_18407(g14817,g12711,g12622);
  nand NAND_18408(g14820,g6307,g12173,g6315,g12423);
  nand NAND_18409(g14822,g12755,g12632);
  nand NAND_18410(g14825,g12806,g12680);
  nand NAND_18411(g14829,g6621,g12137,g6675,g12471);
  nand NAND_18412(g14830,g6605,g12211,g6723,g12721);
  nand NAND_18413(g14838,g12492,g12405);
  nand NAND_18414(g14841,g12593,g12443);
  nand NAND_18415(g14845,g12558,g12798);
  nand NAND_18416(g14848,g12651,g12453);
  nand NAND_18417(g14851,g7738,g12505);
  nand NAND_18418(g14854,g5555,g12093,g5654,g12563);
  nand NAND_18419(g14855,g12700,g12824);
  nand NAND_18420(g14858,g7766,g12515);
  nand NAND_18421(g14861,g12744,g10341);
  nand NAND_18422(g14864,g7791,g10421);
  nand NAND_18423(g14868,g12755,g12680);
  nand NAND_18424(g14871,g6653,g12211,g6661,g12471);
  nand NAND_18425(g14876,g12492,g12443);
  nand NAND_18426(g14879,g12646,g10266);
  nand NAND_18427(g14882,g12558,g12453);
  nand NAND_18428(g14885,g12651,g12505);
  nand NAND_18429(g14889,g12609,g12824);
  nand NAND_18430(g14892,g12700,g12515);
  nand NAND_18431(g14895,g7766,g12571);
  nand NAND_18432(g14898,g5901,g12129,g6000,g12614);
  nand NAND_18433(g14899,g12744,g10421);
  nand NAND_18434(g14902,g7791,g12581);
  nand NAND_18435(g14905,g12785,g7142);
  nand NAND_18436(g14908,g7812,g10491);
  nand NAND_18437(g14915,g12553,g10266);
  nand NAND_18438(g14918,g12646,g12772);
  nand NAND_18439(g14921,g12492,g10266);
  nand NAND_18440(g14924,g12558,g12505);
  nand NAND_18441(g14927,g12695,g10281);
  nand NAND_18442(g14930,g12609,g12515);
  nand NAND_18443(g14933,g12700,g12571);
  nand NAND_18444(g14937,g12667,g10421);
  nand NAND_18445(g14940,g12744,g12581);
  nand NAND_18446(g14943,g7791,g12622);
  nand NAND_18447(g14946,g6247,g12173,g6346,g12672);
  nand NAND_18448(g14947,g12785,g10491);
  nand NAND_18449(g14950,g7812,g12632);
  nand NAND_18450(g14953,g12646,g12405);
  nand NAND_18451(g14956,g12604,g10281);
  nand NAND_18452(g14959,g12695,g12798);
  nand NAND_18453(g14962,g12558,g10281);
  nand NAND_18454(g14965,g12609,g12571);
  nand NAND_18455(g14968,g12739,g10312);
  nand NAND_18456(g14971,g12667,g12581);
  nand NAND_18457(g14974,g12744,g12622);
  nand NAND_18458(g14978,g12716,g10491);
  nand NAND_18459(g14981,g12785,g12632);
  nand NAND_18460(g14984,g7812,g12680);
  nand NAND_18461(g14987,g6593,g12211,g6692,g12721);
  nand NAND_18462(g14993,g12695,g12453);
  nand NAND_18463(g14996,g12662,g10312);
  nand NAND_18464(g14999,g12739,g12824);
  nand NAND_18465(g15002,g12609,g10312);
  nand NAND_18466(g15005,g12667,g12622);
  nand NAND_18467(g15008,g12780,g10341);
  nand NAND_18468(g15011,g12716,g12632);
  nand NAND_18469(g15014,g12785,g12680);
  nand NAND_18470(g15018,g12739,g12515);
  nand NAND_18471(g15021,g12711,g10341);
  nand NAND_18472(g15024,g12780,g10421);
  nand NAND_18473(g15027,g12667,g10341);
  nand NAND_18474(g15030,g12716,g12680);
  nand NAND_18475(g15033,g12806,g7142);
  nand NAND_18476(g15036,g12780,g12581);
  nand NAND_18477(g15039,g12755,g7142);
  nand NAND_18478(g15042,g12806,g10491);
  nand NAND_18479(g15045,g12716,g7142);
  nand NAND_18480(g15572,g12969,g7219);
  nand NAND_18481(g15581,g7232,g12999);
  nand NAND_18482(g15591,g4332,g4322,g13202);
  nand NAND_18483(g15674,g921,g13110);
  nand NAND_18484(g15695,g1266,g13125);
  nand NAND_18485(g15702,g13066,g7293);
  nand NAND_18486(g15708,g7340,g13083);
  nand NAND_18487(g15709,g5224,g14399,g5327,g9780);
  nand NAND_18488(g15710,g319,g13385);
  nand NAND_18489(g15713,g5571,g14425,g5673,g9864);
  nand NAND_18490(g15715,g336,g305,g13385);
  nand NAND_18491(g15717,g10754,g13092);
  nand NAND_18492(g15719,g5256,g14490,g5335,g9780);
  nand NAND_18493(g15720,g5917,g14497,g6019,g9935);
  nand NAND_18494(g15721,g7564,g311,g13385);
  nand NAND_18495(g15723,g10775,g13104);
  nand NAND_18496(g15725,g5603,g14522,g5681,g9864);
  nand NAND_18497(g15726,g6263,g14529,g6365,g10003);
  nand NAND_18498(g15728,g5200,g14399,g5313,g9780);
  nand NAND_18499(g15729,g5949,g14549,g6027,g9935);
  nand NAND_18500(g15730,g6609,g14556,g6711,g10061);
  nand NAND_18501(g15734,g5228,g12059,g5290,g14631);
  nand NAND_18502(g15735,g5547,g14425,g5659,g9864);
  nand NAND_18503(g15736,g6295,g14575,g6373,g10003);
  nand NAND_18504(g15737,g13240,g13115,g7903,g13210);
  nand NAND_18505(g15741,g5244,g14490,g5320,g14631);
  nand NAND_18506(g15742,g5575,g12093,g5637,g14669);
  nand NAND_18507(g15743,g5893,g14497,g6005,g9935);
  nand NAND_18508(g15744,g6641,g14602,g6719,g10061);
  nand NAND_18509(g15748,g13257,g13130,g7922,g13241);
  nand NAND_18510(g15751,g5591,g14522,g5666,g14669);
  nand NAND_18511(g15752,g5921,g12129,g5983,g14701);
  nand NAND_18512(g15753,g6239,g14529,g6351,g10003);
  nand NAND_18513(g15780,g5937,g14549,g6012,g14701);
  nand NAND_18514(g15781,g6267,g12173,g6329,g14745);
  nand NAND_18515(g15782,g6585,g14556,g6697,g10061);
  nand NAND_18516(g15787,g6283,g14575,g6358,g14745);
  nand NAND_18517(g15788,g6613,g12211,g6675,g14786);
  nand NAND_18518(g15798,g6629,g14602,g6704,g14786);
  nand NAND_18519(g15829,g4112,g13831);
  nand NAND_18520(g15832,g7903,g7479,g13256);
  nand NAND_18521(g15833,g14714,g12378,g12337);
  nand NAND_18522(g15843,g7922,g7503,g13264);
  nand NAND_18523(g15844,g14714,g9340,g12378);
  nand NAND_18524(g15853,g14714,g9417,g12337);
  nand NAND_18525(g15864,g14833,g12543,g12487);
  nand NAND_18526(g15867,g14714,g9417,g9340);
  nand NAND_18527(g15877,g14833,g9340,g12543);
  nand NAND_18528(I17379,g13336,g1129);
  nand NAND_18529(I17380,g13336,I17379);
  nand NAND_18530(I17381,g1129,I17379);
  nand NAND_18531(g15904,I17380,I17381);
  nand NAND_18532(g15907,g14833,g9417,g12487);
  nand NAND_18533(I17404,g13378,g1472);
  nand NAND_18534(I17405,g13378,I17404);
  nand NAND_18535(I17406,g1472,I17404);
  nand NAND_18536(g15959,I17405,I17406);
  nand NAND_18537(g15962,g14833,g9417,g9340);
  nand NAND_18538(I17446,g13336,g956);
  nand NAND_18539(I17447,g13336,I17446);
  nand NAND_18540(I17448,g956,I17446);
  nand NAND_18541(g16069,I17447,I17448);
  nand NAND_18542(I17460,g13378,g1300);
  nand NAND_18543(I17461,g13378,I17460);
  nand NAND_18544(I17462,g1300,I17460);
  nand NAND_18545(g16093,I17461,I17462);
  nand NAND_18546(g16097,g13319,g10998);
  nand NAND_18547(I17474,g13336,g1105);
  nand NAND_18548(I17475,g13336,I17474);
  nand NAND_18549(I17476,g1105,I17474);
  nand NAND_18550(g16119,I17475,I17476);
  nand NAND_18551(I17494,g13378,g1448);
  nand NAND_18552(I17495,g13378,I17494);
  nand NAND_18553(I17496,g1448,I17494);
  nand NAND_18554(g16155,I17495,I17496);
  nand NAND_18555(g16181,g13475,g13495,g13057,g13459);
  nand NAND_18556(g16196,g13496,g13513,g13079,g13476);
  nand NAND_18557(g16225,g13544,g13528,g13043);
  nand NAND_18558(g16236,g13573,g13554,g13058);
  nand NAND_18559(g16238,g4698,g13883,g12054);
  nand NAND_18560(g16259,g4743,g13908,g12054);
  nand NAND_18561(g16260,g4888,g13910,g12088);
  nand NAND_18562(g16264,g518,g9158,g13223);
  nand NAND_18563(g16275,g9291,g13480);
  nand NAND_18564(g16278,g8102,g8057,g13664);
  nand NAND_18565(g16281,g4754,g13937,g12054);
  nand NAND_18566(g16282,g4933,g13939,g12088);
  nand NAND_18567(g16291,g13551,g13545);
  nand NAND_18568(g16296,g9360,g13501);
  nand NAND_18569(g16299,g8160,g8112,g13706);
  nand NAND_18570(g16304,g4765,g13970,g12054);
  nand NAND_18571(g16306,g4944,g13971,g12088);
  nand NAND_18572(g16312,g13580,g13574);
  nand NAND_18573(g16316,g9429,g13518);
  nand NAND_18574(g16319,g8224,g8170,g13736);
  nand NAND_18575(g16321,g4955,g13996,g12088);
  nand NAND_18576(g16507,g13797,g13764);
  nand NAND_18577(g16524,g13822,g13798);
  nand NAND_18578(g16586,g13851,g13823);
  nand NAND_18579(g16604,g3251,g11194,g3267,g13877);
  nand NAND_18580(g16625,g3203,g13700,g3274,g11519);
  nand NAND_18581(g16628,g3602,g11207,g3618,g13902);
  nand NAND_18582(g16657,g3554,g13730,g3625,g11576);
  nand NAND_18583(g16660,g3953,g11225,g3969,g13933);
  nand NAND_18584(g16663,g13854,g13834,g14655,g12292);
  nand NAND_18585(I17883,g13336,g1135);
  nand NAND_18586(I17884,g13336,I17883);
  nand NAND_18587(I17885,g1135,I17883);
  nand NAND_18588(g16681,I17884,I17885);
  nand NAND_18589(g16687,g3255,g13700,g3325,g11519);
  nand NAND_18590(g16694,g3905,g13772,g3976,g11631);
  nand NAND_18591(g16696,g13871,g13855,g14682,g12340);
  nand NAND_18592(I17923,g13378,g1478);
  nand NAND_18593(I17924,g13378,I17923);
  nand NAND_18594(I17925,g1478,I17923);
  nand NAND_18595(g16713,I17924,I17925);
  nand NAND_18596(g16719,g3243,g13700,g3310,g11350);
  nand NAND_18597(g16723,g3606,g13730,g3676,g11576);
  nand NAND_18598(g16728,g13884,g13870,g14089,g11639);
  nand NAND_18599(g16741,g3207,g13765,g3303,g11519);
  nand NAND_18600(g16745,g3594,g13730,g3661,g11389);
  nand NAND_18601(g16749,g3957,g13772,g4027,g11631);
  nand NAND_18602(g16757,g13911,g13886,g14120,g11675);
  nand NAND_18603(g16770,g3263,g13765,g3274,g8481);
  nand NAND_18604(g16772,g3558,g13799,g3654,g11576);
  nand NAND_18605(g16776,g3945,g13772,g4012,g11419);
  nand NAND_18606(g16813,g3614,g13799,g3625,g8542);
  nand NAND_18607(g16815,g3909,g13824,g4005,g11631);
  nand NAND_18608(g16854,g3965,g13824,g3976,g8595);
  nand NAND_18609(g16875,g3223,g13765,g3317,g11519);
  nand NAND_18610(g16893,g10685,g13252,g703);
  nand NAND_18611(g16925,g3574,g13799,g3668,g11576);
  nand NAND_18612(g16956,g3925,g13824,g4019,g11631);
  nand NAND_18613(g17137,g13727,g13511,g13527);
  nand NAND_18614(g17217,g7239,g14194);
  nand NAND_18615(g17220,g9369,g9298,g14376);
  nand NAND_18616(g17225,g8612,g14367);
  nand NAND_18617(g17243,g7247,g14212);
  nand NAND_18618(g17246,g9439,g9379,g14405);
  nand NAND_18619(g17287,g7262,g14228);
  nand NAND_18620(g17290,g9506,g9449,g14431);
  nand NAND_18621(g17297,g2729,g14291);
  nand NAND_18622(g17312,g7297,g14248);
  nand NAND_18623(g17315,g9564,g9516,g14503);
  nand NAND_18624(g17363,g8635,g14367);
  nand NAND_18625(g17364,g8639,g14367);
  nand NAND_18626(g17396,g7345,g14272);
  nand NAND_18627(g17399,g9626,g9574,g14535);
  nand NAND_18628(g17412,g14520,g14489);
  nand NAND_18629(g17468,g3215,g13700,g3317,g8481);
  nand NAND_18630(g17474,g14547,g14521);
  nand NAND_18631(g17492,g8655,g14367);
  nand NAND_18632(g17493,g8659,g14367);
  nand NAND_18633(g17495,g3566,g13730,g3668,g8542);
  nand NAND_18634(g17500,g14573,g14548);
  nand NAND_18635(g17513,g3247,g13765,g3325,g8481);
  nand NAND_18636(g17514,g3917,g13772,g4019,g8595);
  nand NAND_18637(g17520,g5260,g12002,g5276,g14631);
  nand NAND_18638(g17525,g14600,g14574);
  nand NAND_18639(I18485,g1677,g14611);
  nand NAND_18640(I18486,g1677,I18485);
  nand NAND_18641(I18487,g14611,I18485);
  nand NAND_18642(g17568,I18486,I18487);
  nand NAND_18643(g17571,g8579,g14367);
  nand NAND_18644(g17572,g3598,g13799,g3676,g8542);
  nand NAND_18645(g17578,g5212,g14399,g5283,g12497);
  nand NAND_18646(g17581,g5607,g12029,g5623,g14669);
  nand NAND_18647(g17586,g14638,g14601);
  nand NAND_18648(I18529,g1811,g14640);
  nand NAND_18649(I18530,g1811,I18529);
  nand NAND_18650(I18531,g14640,I18529);
  nand NAND_18651(g17592,I18530,I18531);
  nand NAND_18652(I18536,g2236,g14642);
  nand NAND_18653(I18537,g2236,I18536);
  nand NAND_18654(I18538,g14642,I18536);
  nand NAND_18655(g17593,I18537,I18538);
  nand NAND_18656(g17595,g8616,g14367);
  nand NAND_18657(g17596,g8686,g14367);
  nand NAND_18658(g17597,g3191,g13700,g3303,g8481);
  nand NAND_18659(g17598,g3949,g13824,g4027,g8595);
  nand NAND_18660(g17605,g5559,g14425,g5630,g12563);
  nand NAND_18661(g17608,g5953,g12067,g5969,g14701);
  nand NAND_18662(I18579,g1945,g14678);
  nand NAND_18663(I18580,g1945,I18579);
  nand NAND_18664(I18581,g14678,I18579);
  nand NAND_18665(g17618,I18580,I18581);
  nand NAND_18666(I18587,g2370,g14679);
  nand NAND_18667(I18588,g2370,I18587);
  nand NAND_18668(I18589,g14679,I18587);
  nand NAND_18669(g17624,I18588,I18589);
  nand NAND_18670(g17634,g3219,g11217,g3281,g13877);
  nand NAND_18671(g17635,g3542,g13730,g3654,g8542);
  nand NAND_18672(g17640,g5264,g14399,g5335,g12497);
  nand NAND_18673(g17647,g5905,g14497,g5976,g12614);
  nand NAND_18674(g17650,g6299,g12101,g6315,g14745);
  nand NAND_18675(I18625,g2079,g14712);
  nand NAND_18676(I18626,g2079,I18625);
  nand NAND_18677(I18627,g14712,I18625);
  nand NAND_18678(g17656,I18626,I18627);
  nand NAND_18679(I18633,g2504,g14713);
  nand NAND_18680(I18634,g2504,I18633);
  nand NAND_18681(I18635,g14713,I18633);
  nand NAND_18682(g17662,I18634,I18635);
  nand NAND_18683(g17668,g3235,g13765,g3310,g13877);
  nand NAND_18684(g17669,g3570,g11238,g3632,g13902);
  nand NAND_18685(g17670,g3893,g13772,g4005,g8595);
  nand NAND_18686(g17675,g5252,g14399,g5320,g12239);
  nand NAND_18687(g17679,g5611,g14425,g5681,g12563);
  nand NAND_18688(g17686,g6251,g14529,g6322,g12672);
  nand NAND_18689(g17689,g6645,g12137,g6661,g14786);
  nand NAND_18690(I18680,g2638,g14752);
  nand NAND_18691(I18681,g2638,I18680);
  nand NAND_18692(I18682,g14752,I18680);
  nand NAND_18693(g17699,I18681,I18682);
  nand NAND_18694(g17705,g3586,g13799,g3661,g13902);
  nand NAND_18695(g17706,g3921,g11255,g3983,g13933);
  nand NAND_18696(g17708,g5216,g14490,g5313,g12497);
  nand NAND_18697(g17712,g5599,g14425,g5666,g12301);
  nand NAND_18698(g17716,g5957,g14497,g6027,g12614);
  nand NAND_18699(g17723,g6597,g14556,g6668,g12721);
  nand NAND_18700(g17732,g3937,g13824,g4012,g13933);
  nand NAND_18701(g17734,g5272,g14490,g5283,g9780);
  nand NAND_18702(g17736,g5563,g14522,g5659,g12563);
  nand NAND_18703(g17740,g5945,g14497,g6012,g12351);
  nand NAND_18704(g17744,g6303,g14529,g6373,g12672);
  nand NAND_18705(g17748,g562,g14708,g12323);
  nand NAND_18706(g17755,g5619,g14522,g5630,g9864);
  nand NAND_18707(g17757,g5909,g14549,g6005,g12614);
  nand NAND_18708(g17761,g6291,g14529,g6358,g12423);
  nand NAND_18709(g17765,g6649,g14556,g6719,g12721);
  nand NAND_18710(g17773,g5965,g14549,g5976,g9935);
  nand NAND_18711(g17775,g6255,g14575,g6351,g12672);
  nand NAND_18712(g17779,g6637,g14556,g6704,g12471);
  nand NAND_18713(g17788,g5232,g14490,g5327,g12497);
  nand NAND_18714(g17790,g6311,g14575,g6322,g10003);
  nand NAND_18715(g17792,g6601,g14602,g6697,g12721);
  nand NAND_18716(g17814,g5579,g14522,g5673,g12563);
  nand NAND_18717(g17816,g6657,g14602,g6668,g10061);
  nand NAND_18718(g17820,g5925,g14549,g6019,g12614);
  nand NAND_18719(g17846,g6271,g14575,g6365,g12672);
  nand NAND_18720(g17872,g6617,g14602,g6711,g12721);
  nand NAND_18721(g19265,g15721,g15715,g13091,g15710);
  nand NAND_18722(g19335,g15717,g1056);
  nand NAND_18723(g19358,g15723,g1399);
  nand NAND_18724(g19442,g11431,g17794);
  nand NAND_18725(g19450,g11471,g17794);
  nand NAND_18726(g19455,g15969,g10841,g7781);
  nand NAND_18727(g19466,g11562,g17794);
  nand NAND_18728(g19474,g11609,g17794);
  nand NAND_18729(g19483,g15969,g10841,g10922);
  nand NAND_18730(g19495,g15969,g10841,g7781);
  nand NAND_18731(g19506,g4087,g15825);
  nand NAND_18732(g19510,g15969,g10841,g10899);
  nand NAND_18733(g19513,g15969,g10841,g10922);
  nand NAND_18734(g19530,g15829,g10841);
  nand NAND_18735(g19546,g15969,g10841,g10884);
  nand NAND_18736(g19549,g15969,g10841,g10899);
  nand NAND_18737(g19589,g15969,g10841,g10884);
  nand NAND_18738(g19597,g1199,g15995);
  nand NAND_18739(g19611,g1070,g1199,g15995);
  nand NAND_18740(g19614,g1542,g16047);
  nand NAND_18741(g19632,g1413,g1542,g16047);
  nand NAND_18742(I20165,g16246,g990);
  nand NAND_18743(I20166,g16246,I20165);
  nand NAND_18744(I20167,g990,I20165);
  nand NAND_18745(g19764,I20166,I20167);
  nand NAND_18746(I20187,g16272,g1333);
  nand NAND_18747(I20188,g16272,I20187);
  nand NAND_18748(I20189,g1333,I20187);
  nand NAND_18749(g19782,I20188,I20189);
  nand NAND_18750(I20203,g16246,g11147);
  nand NAND_18751(I20204,g16246,I20203);
  nand NAND_18752(I20205,g11147,I20203);
  nand NAND_18753(g19792,I20204,I20205);
  nand NAND_18754(g19795,g13600,g16275);
  nand NAND_18755(I20221,g16272,g11170);
  nand NAND_18756(I20222,g16272,I20221);
  nand NAND_18757(I20223,g11170,I20221);
  nand NAND_18758(g19854,I20222,I20223);
  nand NAND_18759(g19856,g13626,g16278,g8105);
  nand NAND_18760(g19857,g13628,g16296);
  nand NAND_18761(g19874,g13665,g16299,g8163);
  nand NAND_18762(g19875,g13667,g16316);
  nand NAND_18763(g19886,g11403,g17794);
  nand NAND_18764(g19903,g13707,g16319,g8227);
  nand NAND_18765(g19913,g11430,g17794);
  nand NAND_18766(g19916,g3029,g16313);
  nand NAND_18767(g19962,g11470,g17794);
  nand NAND_18768(g19965,g3380,g16424);
  nand NAND_18769(g20007,g11512,g17794);
  nand NAND_18770(g20011,g3731,g16476);
  nand NAND_18771(g20039,g11250,g17794);
  nand NAND_18772(g20055,g11269,g17794);
  nand NAND_18773(g20068,g11293,g17794);
  nand NAND_18774(g20076,g13795,g16521);
  nand NAND_18775(g20081,g11325,g17794);
  nand NAND_18776(g20092,g11373,g17794);
  nand NAND_18777(g20107,g11404,g17794);
  nand NAND_18778(g20111,g17513,g14517,g17468,g14422);
  nand NAND_18779(g20133,g17668,g17634,g17597,g14569);
  nand NAND_18780(g20134,g17572,g14542,g17495,g14452);
  nand NAND_18781(g20150,g17705,g17669,g17635,g14590);
  nand NAND_18782(g20151,g17598,g14570,g17514,g14519);
  nand NAND_18783(g20161,g17732,g17706,g17670,g14625);
  nand NAND_18784(g20163,g16663,g13938);
  nand NAND_18785(g20170,g16741,g13897,g16687,g13866);
  nand NAND_18786(g20172,g16876,g8131);
  nand NAND_18787(g20173,g16696,g13972);
  nand NAND_18788(g20181,g13252,g16846);
  nand NAND_18789(g20184,g16770,g13918,g16719,g13896);
  nand NAND_18790(g20185,g16772,g13928,g16723,g13882);
  nand NAND_18791(g20186,g16926,g8177);
  nand NAND_18792(g20198,g16813,g13958,g16745,g13927);
  nand NAND_18793(g20199,g16815,g13968,g16749,g13907);
  nand NAND_18794(I20460,g17515,g14187);
  nand NAND_18795(I20461,g17515,I20460);
  nand NAND_18796(I20462,g14187,I20460);
  nand NAND_18797(g20200,I20461,I20462);
  nand NAND_18798(I20467,g16663,g16728);
  nand NAND_18799(I20468,g16663,I20467);
  nand NAND_18800(I20469,g16728,I20467);
  nand NAND_18801(g20201,I20468,I20469);
  nand NAND_18802(g20214,g16854,g13993,g16776,g13967);
  nand NAND_18803(I20486,g16696,g16757);
  nand NAND_18804(I20487,g16696,I20486);
  nand NAND_18805(I20488,g16757,I20486);
  nand NAND_18806(g20216,I20487,I20488);
  nand NAND_18807(g20236,g16875,g14014,g16625,g16604);
  nand NAND_18808(g20248,g17056,g14146,g14123);
  nand NAND_18809(g20271,g16925,g14054,g16657,g16628);
  nand NAND_18810(g20371,g16956,g14088,g16694,g16660);
  nand NAND_18811(g20619,g14317,g17217);
  nand NAND_18812(g20644,g14342,g17220,g9372);
  nand NAND_18813(g20645,g14344,g17243);
  nand NAND_18814(g20675,g14377,g17246,g9442);
  nand NAND_18815(g20676,g14379,g17287);
  nand NAND_18816(g20733,g14406,g17290,g9509);
  nand NAND_18817(g20734,g14408,g17312);
  nand NAND_18818(g20783,g14616,g17225);
  nand NAND_18819(g20784,g14616,g17595);
  nand NAND_18820(g20838,g5041,g17284);
  nand NAND_18821(g20870,g14432,g17315,g9567);
  nand NAND_18822(g20871,g14434,g17396);
  nand NAND_18823(g20979,g5385,g17309);
  nand NAND_18824(g21011,g14504,g17399,g9629);
  nand NAND_18825(g21124,g5731,g17393);
  nand NAND_18826(g21186,g14616,g17363);
  nand NAND_18827(g21187,g14616,g17364);
  nand NAND_18828(g21190,g6077,g17420);
  nand NAND_18829(g21253,g6423,g17482);
  nand NAND_18830(g21272,g11268,g17157);
  nand NAND_18831(g21283,g11291,g17157);
  nand NAND_18832(g21287,g14616,g17571);
  nand NAND_18833(g21288,g14616,g17492);
  nand NAND_18834(g21289,g14616,g17493);
  nand NAND_18835(g21294,g11324,g17157);
  nand NAND_18836(g21301,g11371,g17157);
  nand NAND_18837(g21307,g15719,g13067,g15709,g13040);
  nand NAND_18838(g21330,g11401,g17157);
  nand NAND_18839(g21331,g11402,g17157);
  nand NAND_18840(g21334,g14616,g17596);
  nand NAND_18841(g21338,g15741,g15734,g15728,g13097);
  nand NAND_18842(g21339,g15725,g13084,g15713,g13050);
  nand NAND_18843(g21344,g11428,g17157);
  nand NAND_18844(g21345,g11429,g17157);
  nand NAND_18845(g21350,g15751,g15742,g15735,g13108);
  nand NAND_18846(g21351,g15729,g13098,g15720,g13069);
  nand NAND_18847(g21353,g11467,g17157);
  nand NAND_18848(g21354,g11468,g17157);
  nand NAND_18849(g21356,g15780,g15752,g15743,g13118);
  nand NAND_18850(g21357,g15736,g13109,g15726,g13086);
  nand NAND_18851(g21359,g11509,g17157);
  nand NAND_18852(g21360,g11510,g17157);
  nand NAND_18853(g21363,g17708,g14664,g17640,g14598);
  nand NAND_18854(g21364,g15787,g15781,g15753,g13131);
  nand NAND_18855(g21365,g15744,g13119,g15730,g13100);
  nand NAND_18856(g21377,g11560,g17157);
  nand NAND_18857(g21384,g17734,g14686,g17675,g14663);
  nand NAND_18858(g21385,g17736,g14696,g17679,g14636);
  nand NAND_18859(g21386,g15798,g15788,g15782,g13139);
  nand NAND_18860(g21388,g11608,g17157);
  nand NAND_18861(g21401,g17755,g14730,g17712,g14695);
  nand NAND_18862(g21402,g17757,g14740,g17716,g14674);
  nand NAND_18863(g21403,g11652,g17157);
  nand NAND_18864(g21415,g17773,g14771,g17740,g14739);
  nand NAND_18865(g21416,g17775,g14781,g17744,g14706);
  nand NAND_18866(g21417,g11677,g17157);
  nand NAND_18867(g21429,g17788,g14803,g17578,g17520);
  nand NAND_18868(g21432,g17790,g14820,g17761,g14780);
  nand NAND_18869(g21433,g17792,g14830,g17765,g14750);
  nand NAND_18870(g21459,g17814,g14854,g17605,g17581);
  nand NAND_18871(g21462,g17816,g14871,g17779,g14829);
  nand NAND_18872(g21509,g17820,g14898,g17647,g17608);
  nand NAND_18873(g21555,g17846,g14946,g17686,g17650);
  nand NAND_18874(g21603,g17872,g14987,g17723,g17689);
  nand NAND_18875(g22306,g4584,g4616,g13202,g19071);
  nand NAND_18876(g22312,g907,g19063);
  nand NAND_18877(g22325,g1252,g19140);
  nand NAND_18878(g22638,g18957,g2886);
  nand NAND_18879(g22642,g7870,g19560);
  nand NAND_18880(g22643,g20136,g18954);
  nand NAND_18881(g22650,g7888,g19581);
  nand NAND_18882(g22651,g20114,g2873);
  nand NAND_18883(g22661,g20136,g94);
  nand NAND_18884(I21976,g7680,g19620);
  nand NAND_18885(I21977,g7680,I21976);
  nand NAND_18886(I21978,g19620,I21976);
  nand NAND_18887(g22663,I21977,I21978);
  nand NAND_18888(g22666,g18957,g2878);
  nand NAND_18889(g22668,g20219,g2912);
  nand NAND_18890(I21992,g7670,g19638);
  nand NAND_18891(I21993,g7670,I21992);
  nand NAND_18892(I21994,g19638,I21992);
  nand NAND_18893(g22681,I21993,I21994);
  nand NAND_18894(g22687,g19560,g7870);
  nand NAND_18895(g22688,g20219,g2936);
  nand NAND_18896(g22709,g1193,g19611);
  nand NAND_18897(g22711,g19581,g7888);
  nand NAND_18898(g22712,g18957,g2864);
  nand NAND_18899(g22713,g20114,g2890);
  nand NAND_18900(g22715,g20114,g2999);
  nand NAND_18901(g22753,g1536,g19632);
  nand NAND_18902(g22754,g20114,g19376);
  nand NAND_18903(g22755,g20136,g18984);
  nand NAND_18904(g22757,g20114,g7891);
  nand NAND_18905(g22833,g1193,g19560,g10666);
  nand NAND_18906(g22836,g18918,g2852);
  nand NAND_18907(g22837,g20219,g2907);
  nand NAND_18908(g22838,g20219,g2960);
  nand NAND_18909(g22839,g20114,g2988);
  nand NAND_18910(g22850,g1536,g19581,g10699);
  nand NAND_18911(g22852,g18957,g2856);
  nand NAND_18912(g22853,g20219,g2922);
  nand NAND_18913(g22864,g7780,g21156);
  nand NAND_18914(g22874,g18918,g2844);
  nand NAND_18915(g22875,g20516,g2980);
  nand NAND_18916(g22885,g9104,g20154);
  nand NAND_18917(g22902,g18957,g2848);
  nand NAND_18918(g22908,g9104,g20175);
  nand NAND_18919(g22921,g20219,g2950);
  nand NAND_18920(g22940,g18918,g2860);
  nand NAND_18921(g22941,g20219,g2970);
  nand NAND_18922(g22984,g20114,g2868);
  nand NAND_18923(g23010,g20516,g2984);
  nand NAND_18924(g23047,g482,g20000);
  nand NAND_18925(g23067,g20887,g10721);
  nand NAND_18926(g23105,g8097,g19887);
  nand NAND_18927(g23112,g21024,g10733);
  nand NAND_18928(g23132,g8155,g19932);
  nand NAND_18929(g23139,g21163,g10756);
  nand NAND_18930(g23167,g8219,g19981);
  nand NAND_18931(g23195,g20136,g37);
  nand NAND_18932(g23210,g18957,g2882);
  nand NAND_18933(g23266,g18918,g2894);
  nand NAND_18934(g23281,g18957,g2898);
  nand NAND_18935(g23286,g6875,g20887);
  nand NAND_18936(g23309,g6905,g21024);
  nand NAND_18937(g23324,g703,g20181);
  nand NAND_18938(g23342,g6928,g21163);
  nand NAND_18939(g23357,g20201,g11231);
  nand NAND_18940(g23379,g20216,g11248);
  nand NAND_18941(g23428,g13945,g20522);
  nand NAND_18942(I22683,g11893,g21434);
  nand NAND_18943(I22684,g11893,I22683);
  nand NAND_18944(I22685,g21434,I22683);
  nand NAND_18945(g23552,I22684,I22685);
  nand NAND_18946(I22710,g11915,g21434);
  nand NAND_18947(I22711,g11915,I22710);
  nand NAND_18948(I22712,g21434,I22710);
  nand NAND_18949(g23575,I22711,I22712);
  nand NAND_18950(I22717,g11916,g21434);
  nand NAND_18951(I22718,g11916,I22717);
  nand NAND_18952(I22719,g21434,I22717);
  nand NAND_18953(g23576,I22718,I22719);
  nand NAND_18954(g23590,g20682,g11111);
  nand NAND_18955(I22753,g11937,g21434);
  nand NAND_18956(I22754,g11937,I22753);
  nand NAND_18957(I22755,g21434,I22753);
  nand NAND_18958(g23616,I22754,I22755);
  nand NAND_18959(I22760,g11939,g21434);
  nand NAND_18960(I22761,g11939,I22760);
  nand NAND_18961(I22762,g21434,I22760);
  nand NAND_18962(g23617,I22761,I22762);
  nand NAND_18963(g23623,g9364,g20717);
  nand NAND_18964(g23630,g20739,g11123);
  nand NAND_18965(I22792,g11956,g21434);
  nand NAND_18966(I22793,g11956,I22792);
  nand NAND_18967(I22794,g21434,I22792);
  nand NAND_18968(g23655,I22793,I22794);
  nand NAND_18969(I22799,g11960,g21434);
  nand NAND_18970(I22800,g11960,I22799);
  nand NAND_18971(I22801,g21434,I22799);
  nand NAND_18972(g23656,I22800,I22801);
  nand NAND_18973(g23659,g9434,g20854);
  nand NAND_18974(g23666,g20875,g11139);
  nand NAND_18975(I22822,g11978,g21434);
  nand NAND_18976(I22823,g11978,I22822);
  nand NAND_18977(I22824,g21434,I22822);
  nand NAND_18978(g23685,I22823,I22824);
  nand NAND_18979(g23692,g9501,g20995);
  nand NAND_18980(g23699,g21012,g11160);
  nand NAND_18981(I22844,g12113,g21228);
  nand NAND_18982(I22845,g12113,I22844);
  nand NAND_18983(I22846,g21228,I22844);
  nand NAND_18984(g23719,I22845,I22846);
  nand NAND_18985(g23726,g9559,g21140);
  nand NAND_18986(g23733,g20751,g11178);
  nand NAND_18987(I22864,g12146,g21228);
  nand NAND_18988(I22865,g12146,I22864);
  nand NAND_18989(I22866,g21228,I22864);
  nand NAND_18990(g23747,I22865,I22866);
  nand NAND_18991(I22871,g12150,g21228);
  nand NAND_18992(I22872,g12150,I22871);
  nand NAND_18993(I22873,g21228,I22871);
  nand NAND_18994(g23748,I22872,I22873);
  nand NAND_18995(g23756,g9621,g21206);
  nand NAND_18996(I22892,g12189,g21228);
  nand NAND_18997(I22893,g12189,I22892);
  nand NAND_18998(I22894,g21228,I22892);
  nand NAND_18999(g23761,I22893,I22894);
  nand NAND_19000(I22899,g12193,g21228);
  nand NAND_19001(I22900,g12193,I22899);
  nand NAND_19002(I22901,g21228,I22899);
  nand NAND_19003(g23762,I22900,I22901);
  nand NAND_19004(I22921,g14677,g21284);
  nand NAND_19005(I22922,g14677,I22921);
  nand NAND_19006(I22923,g21284,I22921);
  nand NAND_19007(g23778,I22922,I22923);
  nand NAND_19008(I22929,g12223,g21228);
  nand NAND_19009(I22930,g12223,I22929);
  nand NAND_19010(I22931,g21228,I22929);
  nand NAND_19011(g23780,I22930,I22931);
  nand NAND_19012(I22936,g12226,g21228);
  nand NAND_19013(I22937,g12226,I22936);
  nand NAND_19014(I22938,g21228,I22936);
  nand NAND_19015(g23781,I22937,I22938);
  nand NAND_19016(g23782,g2741,g21062);
  nand NAND_19017(I22944,g9492,g19620);
  nand NAND_19018(I22945,g9492,I22944);
  nand NAND_19019(I22946,g19620,I22944);
  nand NAND_19020(g23786,I22945,I22946);
  nand NAND_19021(I22965,g12288,g21228);
  nand NAND_19022(I22966,g12288,I22965);
  nand NAND_19023(I22967,g21228,I22965);
  nand NAND_19024(g23809,I22966,I22967);
  nand NAND_19025(I22972,g9657,g19638);
  nand NAND_19026(I22973,g9657,I22972);
  nand NAND_19027(I22974,g19638,I22972);
  nand NAND_19028(g23810,I22973,I22974);
  nand NAND_19029(g23850,g12185,g19462);
  nand NAND_19030(g23890,g7004,g20682);
  nand NAND_19031(g23909,g7028,g20739);
  nand NAND_19032(g23932,g7051,g20875);
  nand NAND_19033(g23949,g7074,g21012);
  nand NAND_19034(g23972,g7097,g20751);
  nand NAND_19035(I23118,g20076,g417);
  nand NAND_19036(I23119,g20076,I23118);
  nand NAND_19037(I23120,g417,I23118);
  nand NAND_19038(g23975,I23119,I23120);
  nand NAND_19039(g23978,g572,g21389,g12323);
  nand NAND_19040(g24362,g21370,g22136);
  nand NAND_19041(I23585,g22409,g4332);
  nand NAND_19042(I23586,g22409,I23585);
  nand NAND_19043(I23587,g4332,I23585);
  nand NAND_19044(g24369,I23586,I23587);
  nand NAND_19045(I23600,g22360,g4322);
  nand NAND_19046(I23601,g22360,I23600);
  nand NAND_19047(I23602,g4322,I23600);
  nand NAND_19048(g24380,I23601,I23602);
  nand NAND_19049(g24528,g4098,g22654);
  nand NAND_19050(g24544,g22666,g22661,g22651);
  nand NAND_19051(g24547,g22638,g22643,g22754);
  nand NAND_19052(g24566,g22755,g22713);
  nand NAND_19053(g24567,g22957,g2917);
  nand NAND_19054(g24570,g22957,g2941);
  nand NAND_19055(g24574,g22709,g22687);
  nand NAND_19056(g24576,g22957,g2902);
  nand NAND_19057(g24583,g22753,g22711);
  nand NAND_19058(g24584,g22852,g22836,g22715);
  nand NAND_19059(g24591,g22833,g22642);
  nand NAND_19060(g24601,g22957,g2965);
  nand NAND_19061(g24609,g22850,g22650);
  nand NAND_19062(g24620,g22902,g22874);
  nand NAND_19063(g24621,g22957,g2927);
  nand NAND_19064(g24652,g22712,g22940,g22757);
  nand NAND_19065(g24661,g23210,g23195,g22984);
  nand NAND_19066(g24662,g22957,g2955);
  nand NAND_19067(g24677,g22957,g2975);
  nand NAND_19068(g24678,g22994,g23010);
  nand NAND_19069(I23917,g23975,g9333);
  nand NAND_19070(I23918,g23975,I23917);
  nand NAND_19071(I23919,g9333,I23917);
  nand NAND_19072(g24760,I23918,I23919);
  nand NAND_19073(g24776,g3040,g23052);
  nand NAND_19074(g24787,g3391,g23079);
  nand NAND_19075(I23949,g23162,g13603);
  nand NAND_19076(I23950,g23162,I23949);
  nand NAND_19077(I23951,g13603,I23949);
  nand NAND_19078(g24792,I23950,I23951);
  nand NAND_19079(g24793,g3742,g23124);
  nand NAND_19080(I23961,g23184,g13631);
  nand NAND_19081(I23962,g23184,I23961);
  nand NAND_19082(I23963,g13631,I23961);
  nand NAND_19083(g24798,I23962,I23963);
  nand NAND_19084(I23969,g22202,g490);
  nand NAND_19085(I23970,g22202,I23969);
  nand NAND_19086(I23971,g490,I23969);
  nand NAND_19087(g24802,I23970,I23971);
  nand NAND_19088(g24804,g19916,g23105);
  nand NAND_19089(I23978,g23198,g13670);
  nand NAND_19090(I23979,g23198,I23978);
  nand NAND_19091(I23980,g13670,I23978);
  nand NAND_19092(g24807,I23979,I23980);
  nand NAND_19093(I23985,g22182,g482);
  nand NAND_19094(I23986,g22182,I23985);
  nand NAND_19095(I23987,g482,I23985);
  nand NAND_19096(g24808,I23986,I23987);
  nand NAND_19097(g24809,g19965,g23132);
  nand NAND_19098(g24814,g20011,g23167);
  nand NAND_19099(g24880,g23281,g23266,g22839);
  nand NAND_19100(g24890,g13852,g22929);
  nand NAND_19101(g24905,g534,g23088);
  nand NAND_19102(g24906,g8743,g23088);
  nand NAND_19103(g24916,g19450,g23154);
  nand NAND_19104(g24917,g19913,g23172);
  nand NAND_19105(g24918,g136,g23088);
  nand NAND_19106(g24924,g20007,g23172);
  nand NAND_19107(g24925,g20092,g23154);
  nand NAND_19108(g24926,g20172,g20163,g23357,g13995);
  nand NAND_19109(g24932,g19886,g23172);
  nand NAND_19110(g24933,g19466,g23154);
  nand NAND_19111(g24934,g21283,g23462);
  nand NAND_19112(g24936,g20186,g20173,g23379,g14029);
  nand NAND_19113(g24942,g20039,g23172);
  nand NAND_19114(g24943,g20068,g23172);
  nand NAND_19115(g24944,g21354,g23363);
  nand NAND_19116(g24950,g19442,g23154);
  nand NAND_19117(g24951,g199,g23088);
  nand NAND_19118(g24957,g21359,g23462);
  nand NAND_19119(g24958,g21330,g23462);
  nand NAND_19120(g24972,g19962,g23172);
  nand NAND_19121(g24973,g21272,g23462);
  nand NAND_19122(g24974,g21301,g23363);
  nand NAND_19123(g24975,g21388,g23363);
  nand NAND_19124(g24988,g546,g23088);
  nand NAND_19125(g24989,g21345,g23363);
  nand NAND_19126(g25002,g19474,g23154);
  nand NAND_19127(g25003,g21353,g23462);
  nand NAND_19128(g25018,g20107,g23154);
  nand NAND_19129(g25019,g20055,g23172);
  nand NAND_19130(g25020,g21377,g23462);
  nand NAND_19131(g25021,g21417,g23363);
  nand NAND_19132(g25038,g21331,g23363);
  nand NAND_19133(g25048,g542,g23088);
  nand NAND_19134(g25049,g21344,g23462);
  nand NAND_19135(g25062,g21403,g23363);
  nand NAND_19136(g25172,g5052,g23560);
  nand NAND_19137(g25186,g5396,g23602);
  nand NAND_19138(I24363,g23687,g14320);
  nand NAND_19139(I24364,g23687,I24363);
  nand NAND_19140(I24365,g14320,I24363);
  nand NAND_19141(g25199,I24364,I24365);
  nand NAND_19142(g25200,g5742,g23642);
  nand NAND_19143(I24383,g23721,g14347);
  nand NAND_19144(I24384,g23721,I24383);
  nand NAND_19145(I24385,g14347,I24383);
  nand NAND_19146(g25215,I24384,I24385);
  nand NAND_19147(g25216,g6088,g23678);
  nand NAND_19148(g25233,g20838,g23623);
  nand NAND_19149(I24414,g23751,g14382);
  nand NAND_19150(I24415,g23751,I24414);
  nand NAND_19151(I24416,g14382,I24414);
  nand NAND_19152(g25236,I24415,I24416);
  nand NAND_19153(g25237,g6434,g23711);
  nand NAND_19154(g25255,g20979,g23659);
  nand NAND_19155(I24438,g23771,g14411);
  nand NAND_19156(I24439,g23771,I24438);
  nand NAND_19157(I24440,g14411,I24438);
  nand NAND_19158(g25258,I24439,I24440);
  nand NAND_19159(g25268,g21124,g23692);
  nand NAND_19160(I24461,g23796,g14437);
  nand NAND_19161(I24462,g23796,I24461);
  nand NAND_19162(I24463,g14437,I24461);
  nand NAND_19163(g25271,I24462,I24463);
  nand NAND_19164(g25275,g22342,g11991);
  nand NAND_19165(g25293,g21190,g23726);
  nand NAND_19166(g25300,g22369,g12018);
  nand NAND_19167(g25309,g22384,g12021);
  nand NAND_19168(g25334,g21253,g23756);
  nand NAND_19169(g25337,g22342,g1648,g8187);
  nand NAND_19170(g25341,g22417,g12047);
  nand NAND_19171(g25349,g22432,g12051);
  nand NAND_19172(g25381,g538,g23088);
  nand NAND_19173(g25382,g12333,g22342);
  nand NAND_19174(g25385,g22369,g1783,g8241);
  nand NAND_19175(g25389,g22457,g12082);
  nand NAND_19176(g25396,g22384,g2208,g8259);
  nand NAND_19177(g25400,g22472,g12086);
  nand NAND_19178(g25425,g20081,g23172);
  nand NAND_19179(g25426,g12371,g22369);
  nand NAND_19180(g25429,g22417,g1917,g8302);
  nand NAND_19181(g25432,g12374,g22384);
  nand NAND_19182(g25435,g22432,g2342,g8316);
  nand NAND_19183(g25439,g22498,g12122);
  nand NAND_19184(g25467,g12432,g22417);
  nand NAND_19185(g25470,g22457,g2051,g8365);
  nand NAND_19186(g25473,g12437,g22432);
  nand NAND_19187(g25476,g22472,g2476,g8373);
  nand NAND_19188(g25492,g12479,g22457);
  nand NAND_19189(g25495,g12483,g22472);
  nand NAND_19190(g25498,g22498,g2610,g8418);
  nand NAND_19191(g25514,g12540,g22498);
  nand NAND_19192(g25527,g21294,g23462);
  nand NAND_19193(g25531,g22763,g2868);
  nand NAND_19194(g25532,g21360,g23363);
  nand NAND_19195(g25537,g22763,g2873);
  nand NAND_19196(g25779,g19694,g24362);
  nand NAND_19197(g25888,g914,g24439);
  nand NAND_19198(g25895,g1259,g24453);
  nand NAND_19199(g25953,g22756,g24570,g22688);
  nand NAND_19200(g25974,g24576,g22837);
  nand NAND_19201(g25984,g24567,g22668);
  nand NAND_19202(g25985,g24631,g23956);
  nand NAND_19203(g25995,g24621,g22853);
  nand NAND_19204(g25996,g24601,g22838);
  nand NAND_19205(g26025,g22405,g24631);
  nand NAND_19206(g26052,g22714,g24662,g22921);
  nand NAND_19207(g26053,g22875,g24677,g22941);
  nand NAND_19208(g26208,g7975,g24751);
  nand NAND_19209(g26235,g8016,g24766);
  nand NAND_19210(I25219,g482,g24718);
  nand NAND_19211(I25220,g482,I25219);
  nand NAND_19212(I25221,g24718,I25219);
  nand NAND_19213(g26248,I25220,I25221);
  nand NAND_19214(g26255,g8075,g24779);
  nand NAND_19215(I25242,g490,g24744);
  nand NAND_19216(I25243,g490,I25242);
  nand NAND_19217(I25244,g24744,I25242);
  nand NAND_19218(g26269,I25243,I25244);
  nand NAND_19219(g26352,g744,g24875,g11679);
  nand NAND_19220(g26382,g577,g24953,g12323);
  nand NAND_19221(g26666,g9229,g25144);
  nand NAND_19222(g26685,g9264,g25160);
  nand NAND_19223(g26714,g9316,g25175);
  nand NAND_19224(g26745,g6856,g25317);
  nand NAND_19225(g26752,g9397,g25189);
  nand NAND_19226(g26782,g9467,g25203);
  nand NAND_19227(I25845,g26212,g24799);
  nand NAND_19228(I25846,g26212,I25845);
  nand NAND_19229(I25847,g24799,I25845);
  nand NAND_19230(g27141,I25846,I25847);
  nand NAND_19231(I25907,g26256,g24782);
  nand NAND_19232(I25908,g26256,I25907);
  nand NAND_19233(I25909,g24782,I25907);
  nand NAND_19234(g27223,I25908,I25909);
  nand NAND_19235(g27273,g10504,g26131,g26105);
  nand NAND_19236(g27282,g11192,g26269,g26248,g479);
  nand NAND_19237(g27295,g24776,g26208);
  nand NAND_19238(g27306,g24787,g26235);
  nand NAND_19239(g27317,g24793,g26255);
  nand NAND_19240(I26049,g25997,g13500);
  nand NAND_19241(I26050,g25997,I26049);
  nand NAND_19242(I26051,g13500,I26049);
  nand NAND_19243(g27365,I26050,I26051);
  nand NAND_19244(g27377,g10685,g25930);
  nand NAND_19245(I26070,g26026,g13517);
  nand NAND_19246(I26071,g26026,I26070);
  nand NAND_19247(I26072,g13517,I26070);
  nand NAND_19248(g27380,I26071,I26072);
  nand NAND_19249(I26093,g26055,g13539);
  nand NAND_19250(I26094,g26055,I26093);
  nand NAND_19251(I26095,g13539,I26093);
  nand NAND_19252(g27401,I26094,I26095);
  nand NAND_19253(g27463,g287,g26330,g23204);
  nand NAND_19254(g27468,g24951,g24932,g24925,g26852);
  nand NAND_19255(g27550,g24943,g25772);
  nand NAND_19256(g27577,g25019,g25002,g24988,g25765);
  nand NAND_19257(g27582,g10857,g26131,g26105);
  nand NAND_19258(g27586,g24924,g24916,g24905,g26863);
  nand NAND_19259(g27587,g24917,g25018,g24918,g26857);
  nand NAND_19260(g27593,g24972,g24950,g24906,g26861);
  nand NAND_19261(g27613,g24942,g24933,g25048,g26871);
  nand NAND_19262(g27654,g164,g26598,g23042);
  nand NAND_19263(g27670,g25172,g26666);
  nand NAND_19264(g27679,g25186,g26685);
  nand NAND_19265(g27687,g25200,g26714);
  nand NAND_19266(g27693,g25216,g26752);
  nand NAND_19267(g27705,g25237,g26782);
  nand NAND_19268(g27738,g21228,g25243,g26424,g26148);
  nand NAND_19269(I26366,g26400,g14211);
  nand NAND_19270(I26367,g26400,I26366);
  nand NAND_19271(I26368,g14211,I26366);
  nand NAND_19272(g27767,I26367,I26368);
  nand NAND_19273(g27775,g21228,g25262,g26424,g26166);
  nand NAND_19274(g27796,g21228,g25263,g26424,g26171);
  nand NAND_19275(I26393,g26488,g14227);
  nand NAND_19276(I26394,g26488,I26393);
  nand NAND_19277(I26395,g14227,I26393);
  nand NAND_19278(g27824,I26394,I26395);
  nand NAND_19279(g27833,g21228,g25282,g26424,g26190);
  nand NAND_19280(g27854,g21228,g25283,g26424,g26195);
  nand NAND_19281(I26417,g26519,g14247);
  nand NAND_19282(I26418,g26519,I26417);
  nand NAND_19283(I26419,g14247,I26417);
  nand NAND_19284(g27876,I26418,I26419);
  nand NAND_19285(g27882,g21228,g25307,g26424,g26213);
  nand NAND_19286(g27903,g21228,g25316,g26424,g26218);
  nand NAND_19287(I26438,g26549,g14271);
  nand NAND_19288(I26439,g26549,I26438);
  nand NAND_19289(I26440,g14271,I26438);
  nand NAND_19290(g27925,I26439,I26440);
  nand NAND_19291(g27931,g25425,g25381,g25780);
  nand NAND_19292(g27933,g21228,g25356,g26424,g26236);
  nand NAND_19293(I26459,g26576,g14306);
  nand NAND_19294(I26460,g26576,I26459);
  nand NAND_19295(I26461,g14306,I26459);
  nand NAND_19296(g27955,I26460,I26461);
  nand NAND_19297(g28109,g27051,g25783);
  nand NAND_19298(g28131,g27051,g25838);
  nand NAND_19299(g28167,g925,g27046);
  nand NAND_19300(g28174,g1270,g27059);
  nand NAND_19301(g28203,g12546,g27985,g27977);
  nand NAND_19302(g28206,g12546,g26105,g27985);
  nand NAND_19303(g28207,g12546,g26131,g27977);
  nand NAND_19304(g28259,g10504,g26987,g26973);
  nand NAND_19305(g28270,g10504,g26105,g26987);
  nand NAND_19306(g28271,g10533,g27004,g26990);
  nand NAND_19307(g28287,g10504,g26131,g26973);
  nand NAND_19308(g28288,g10533,g26105,g27004);
  nand NAND_19309(g28298,g10533,g26131,g26990);
  nand NAND_19310(g28336,g27064,g24756,g27163,g19644);
  nand NAND_19311(g28349,g27074,g24770,g27187,g19644);
  nand NAND_19312(g28363,g27064,g13593);
  nand NAND_19313(g28376,g27064,g13620);
  nand NAND_19314(g28381,g27074,g13621);
  nand NAND_19315(g28391,g27064,g13637);
  nand NAND_19316(g28395,g27074,g13655);
  nand NAND_19317(g28406,g27064,g13675);
  nand NAND_19318(g28410,g27074,g13679);
  nand NAND_19319(g28421,g27074,g13715);
  nand NAND_19320(g28448,g23975,g27377);
  nand NAND_19321(g28500,g590,g27629,g12323);
  nand NAND_19322(g28504,g758,g27528,g11679);
  nand NAND_19323(g28512,g10857,g27155,g27142);
  nand NAND_19324(g28516,g10857,g26105,g27155);
  nand NAND_19325(g28522,g10857,g26131,g27142);
  nand NAND_19326(g28736,g27742,g7308,g7252);
  nand NAND_19327(g28755,g27742,g7268,g1592);
  nand NAND_19328(g28758,g27779,g7356,g7275);
  nand NAND_19329(g28765,g27800,g7374,g7280);
  nand NAND_19330(g28780,g27742,g7308,g1636);
  nand NAND_19331(g28783,g27779,g7315,g1728);
  nand NAND_19332(g28786,g27837,g7405,g7322);
  nand NAND_19333(g28793,g27800,g7328,g2153);
  nand NAND_19334(g28796,g27858,g7418,g7335);
  nand NAND_19335(g28820,g27742,g1668,g1592);
  nand NAND_19336(g28823,g27738,g14565);
  nand NAND_19337(g28824,g27779,g7356,g1772);
  nand NAND_19338(g28827,g27837,g7362,g1862);
  nand NAND_19339(g28830,g27886,g7451,g7369);
  nand NAND_19340(g28837,g27800,g7374,g2197);
  nand NAND_19341(g28840,g27858,g7380,g2287);
  nand NAND_19342(g28843,g27907,g7456,g7387);
  nand NAND_19343(g28853,g27742,g1636,g7252);
  nand NAND_19344(g28856,g27738,g8093);
  nand NAND_19345(g28857,g27779,g1802,g1728);
  nand NAND_19346(g28860,g27775,g14586);
  nand NAND_19347(g28861,g27837,g7405,g1906);
  nand NAND_19348(g28864,g27886,g7411,g1996);
  nand NAND_19349(g28867,g27800,g2227,g2153);
  nand NAND_19350(g28870,g27796,g14588);
  nand NAND_19351(g28871,g27858,g7418,g2331);
  nand NAND_19352(g28874,g27907,g7424,g2421);
  nand NAND_19353(g28877,g27937,g7490,g7431);
  nand NAND_19354(g28885,g27742,g1668,g7268);
  nand NAND_19355(g28888,g27738,g8139);
  nand NAND_19356(g28892,g27779,g1772,g7275);
  nand NAND_19357(g28895,g27775,g8146);
  nand NAND_19358(g28896,g27837,g1936,g1862);
  nand NAND_19359(g28899,g27833,g14612);
  nand NAND_19360(g28900,g27886,g7451,g2040);
  nand NAND_19361(g28903,g27800,g2197,g7280);
  nand NAND_19362(g28906,g27796,g8150);
  nand NAND_19363(g28907,g27858,g2361,g2287);
  nand NAND_19364(g28910,g27854,g14614);
  nand NAND_19365(g28911,g27907,g7456,g2465);
  nand NAND_19366(g28914,g27937,g7462,g2555);
  nand NAND_19367(g28920,g27779,g1802,g7315);
  nand NAND_19368(g28923,g27775,g8195);
  nand NAND_19369(g28927,g27837,g1906,g7322);
  nand NAND_19370(g28930,g27833,g8201);
  nand NAND_19371(g28931,g27886,g2070,g1996);
  nand NAND_19372(g28934,g27882,g14641);
  nand NAND_19373(g28935,g27800,g2227,g7328);
  nand NAND_19374(g28938,g27796,g8205);
  nand NAND_19375(g28942,g27858,g2331,g7335);
  nand NAND_19376(g28945,g27854,g8211);
  nand NAND_19377(g28946,g27907,g2495,g2421);
  nand NAND_19378(g28949,g27903,g14643);
  nand NAND_19379(g28950,g27937,g7490,g2599);
  nand NAND_19380(g28955,g27837,g1936,g7362);
  nand NAND_19381(g28958,g27833,g8249);
  nand NAND_19382(g28962,g27886,g2040,g7369);
  nand NAND_19383(g28965,g27882,g8255);
  nand NAND_19384(g28966,g27858,g2361,g7380);
  nand NAND_19385(g28969,g27854,g8267);
  nand NAND_19386(g28973,g27907,g2465,g7387);
  nand NAND_19387(g28976,g27903,g8273);
  nand NAND_19388(g28977,g27937,g2629,g2555);
  nand NAND_19389(g28980,g27933,g14680);
  nand NAND_19390(g28987,g27886,g2070,g7411);
  nand NAND_19391(g28990,g27882,g8310);
  nand NAND_19392(g28994,g27907,g2495,g7424);
  nand NAND_19393(g28997,g27903,g8324);
  nand NAND_19394(g29001,g27937,g2599,g7431);
  nand NAND_19395(g29004,g27933,g8330);
  nand NAND_19396(g29015,g27742,g9586);
  nand NAND_19397(g29018,g9586,g27742);
  nand NAND_19398(g29025,g27937,g2629,g7462);
  nand NAND_19399(g29028,g27933,g8381);
  nand NAND_19400(g29046,g27779,g9640);
  nand NAND_19401(g29049,g9640,g27779);
  nand NAND_19402(g29057,g27800,g9649);
  nand NAND_19403(g29060,g9649,g27800);
  nand NAND_19404(g29082,g27837,g9694);
  nand NAND_19405(g29085,g9694,g27837);
  nand NAND_19406(g29094,g27858,g9700);
  nand NAND_19407(g29097,g9700,g27858);
  nand NAND_19408(g29118,g27886,g9755);
  nand NAND_19409(g29121,g9755,g27886);
  nand NAND_19410(g29131,g27907,g9762);
  nand NAND_19411(g29134,g9762,g27907);
  nand NAND_19412(g29154,g27937,g9835);
  nand NAND_19413(g29157,g9835,g27937);
  nand NAND_19414(g29186,g27051,g4507);
  nand NAND_19415(g29335,g25540,g28131);
  nand NAND_19416(g29355,g24383,g28109);
  nand NAND_19417(g29540,g28336,g13464);
  nand NAND_19418(g29556,g28349,g13486);
  nand NAND_19419(g29657,g28363,g13634);
  nand NAND_19420(g29660,g28448,g9582);
  nand NAND_19421(g29672,g28376,g13672);
  nand NAND_19422(g29676,g28381,g13676);
  nand NAND_19423(g29679,g153,g28353,g23042);
  nand NAND_19424(g29694,g28391,g13709);
  nand NAND_19425(g29702,g28395,g13712);
  nand NAND_19426(g29719,g28406,g13739);
  nand NAND_19427(g29722,g28410,g13742);
  nand NAND_19428(g29737,g28421,g13779);
  nand NAND_19429(g29778,g294,g28444,g23204);
  nand NAND_19430(g30573,g29355,g19666);
  nand NAND_19431(g30580,g29335,g19666);
  nand NAND_19432(g31003,g27163,g29497,g19644);
  nand NAND_19433(g31009,g27187,g29503,g19644);
  nand NAND_19434(g31262,g767,g29916,g11679);
  nand NAND_19435(g31509,g599,g29933,g12323);
  nand NAND_19436(I29253,g29482,g12017);
  nand NAND_19437(I29254,g29482,I29253);
  nand NAND_19438(I29255,g12017,I29253);
  nand NAND_19439(g31669,I29254,I29255);
  nand NAND_19440(I29261,g29485,g12046);
  nand NAND_19441(I29262,g29485,I29261);
  nand NAND_19442(I29263,g12046,I29261);
  nand NAND_19443(g31671,I29262,I29263);
  nand NAND_19444(I29269,g29486,g12050);
  nand NAND_19445(I29270,g29486,I29269);
  nand NAND_19446(I29271,g12050,I29269);
  nand NAND_19447(g31706,I29270,I29271);
  nand NAND_19448(I29277,g29488,g12081);
  nand NAND_19449(I29278,g29488,I29277);
  nand NAND_19450(I29279,g12081,I29277);
  nand NAND_19451(g31708,I29278,I29279);
  nand NAND_19452(I29284,g29489,g12085);
  nand NAND_19453(I29285,g29489,I29284);
  nand NAND_19454(I29286,g12085,I29284);
  nand NAND_19455(g31709,I29285,I29286);
  nand NAND_19456(I29295,g29495,g12117);
  nand NAND_19457(I29296,g29495,I29295);
  nand NAND_19458(I29297,g12117,I29295);
  nand NAND_19459(g31747,I29296,I29297);
  nand NAND_19460(I29302,g29496,g12121);
  nand NAND_19461(I29303,g29496,I29302);
  nand NAND_19462(I29304,g12121,I29302);
  nand NAND_19463(g31748,I29303,I29304);
  nand NAND_19464(I29313,g29501,g12154);
  nand NAND_19465(I29314,g29501,I29313);
  nand NAND_19466(I29315,g12154,I29313);
  nand NAND_19467(g31753,I29314,I29315);
  nand NAND_19468(g31950,g7285,g30573);
  nand NAND_19469(g31971,g30573,g10511);
  nand NAND_19470(g31978,g30580,g15591);
  nand NAND_19471(g31997,g22306,g30580);
  nand NAND_19472(g32057,g31003,g13297);
  nand NAND_19473(g32072,g31009,g13301);
  nand NAND_19474(g33083,g7805,g32118);
  nand NAND_19475(g33299,g608,g32296,g12323);
  nand NAND_19476(g33306,g776,g32212,g11679);
  nand NAND_19477(g33394,g10159,g4474,g32426);
  nand NAND_19478(g33669,g33378,g862);
  nand NAND_19479(g33679,g33394,g10737,g10308);
  nand NAND_19480(g33838,g33083,g4369);
  nand NAND_19481(g33925,g33394,g4462,g4467);
  nand NAND_19482(g33930,g33394,g12767,g9848);
  nand NAND_19483(g33933,g33394,g12491,g12819,g12796);
  nand NAND_19484(g34048,g33669,g10583,g7442);
  nand NAND_19485(I31972,g33641,g33631);
  nand NAND_19486(I31973,g33641,I31972);
  nand NAND_19487(I31974,g33631,I31972);
  nand NAND_19488(g34051,I31973,I31974);
  nand NAND_19489(I31983,g33653,g33648);
  nand NAND_19490(I31984,g33653,I31983);
  nand NAND_19491(I31985,g33648,I31983);
  nand NAND_19492(g34056,I31984,I31985);
  nand NAND_19493(g34162,g785,g33823,g11679);
  nand NAND_19494(g34174,g617,g33851,g12323);
  nand NAND_19495(I32185,g33665,g33661);
  nand NAND_19496(I32186,g33665,I32185);
  nand NAND_19497(I32187,g33661,I32185);
  nand NAND_19498(g34220,I32186,I32187);
  nand NAND_19499(I32202,g33937,g33670);
  nand NAND_19500(I32203,g33937,I32202);
  nand NAND_19501(I32204,g33670,I32202);
  nand NAND_19502(g34227,I32203,I32204);
  nand NAND_19503(I32431,g34056,g34051);
  nand NAND_19504(I32432,g34056,I32431);
  nand NAND_19505(I32433,g34051,I32431);
  nand NAND_19506(g34422,I32432,I32433);
  nand NAND_19507(I32439,g34227,g34220);
  nand NAND_19508(I32440,g34227,I32439);
  nand NAND_19509(I32441,g34220,I32439);
  nand NAND_19510(g34424,I32440,I32441);
  nand NAND_19511(I32516,g34424,g34422);
  nand NAND_19512(I32517,g34424,I32516);
  nand NAND_19513(I32518,g34422,I32516);
  nand NAND_19514(g34469,I32517,I32518);
  nand NAND_19515(g34545,g11679,g794,g34354);
  nand NAND_19516(g34550,g626,g34359,g12323);
  nand NAND_19517(I32756,g34469,g25779);
  nand NAND_19518(I32757,g34469,I32756);
  nand NAND_19519(I32758,g25779,I32756);
  nand NAND_19520(g34650,I32757,I32758);
  nor NOR_19521(g7139,g5406,g5366);
  nor NOR_19522(g7142,g6573,g6565);
  nor NOR_19523(g7158,g5752,g5712);
  nor NOR_19524(g7175,g6098,g6058);
  nor NOR_19525(g7192,g6444,g6404);
  nor NOR_19526(g7304,g1183,g1171);
  nor NOR_19527(g7352,g1526,g1514);
  nor NOR_19528(g7499,g333,g355);
  nor NOR_19529(g7567,g979,g990);
  nor NOR_19530(g7601,g1322,g1333);
  nor NOR_19531(g7661,g1211,g1216,g1221,g1205);
  nor NOR_19532(g7675,g1554,g1559,g1564,g1548);
  nor NOR_19533(g7781,g4064,g4057);
  nor NOR_19534(g8086,g168,g174,g182);
  nor NOR_19535(g8131,g4776,g4801,g4793);
  nor NOR_19536(g8177,g4966,g4991,g4983);
  nor NOR_19537(g8182,g405,g392);
  nor NOR_19538(g8720,g358,g365);
  nor NOR_19539(g8864,g3179,g3171);
  nor NOR_19540(g8906,g3530,g3522);
  nor NOR_19541(g8933,g4709,g4785);
  nor NOR_19542(g8958,g3881,g3873);
  nor NOR_19543(g8984,g4899,g4975);
  nor NOR_19544(g9015,g3050,g3010);
  nor NOR_19545(g9061,g3401,g3361);
  nor NOR_19546(g9100,g3752,g3712);
  nor NOR_19547(g9586,g1668,g1592);
  nor NOR_19548(g9602,g4688,g4681,g4674,g4646);
  nor NOR_19549(g9640,g1802,g1728);
  nor NOR_19550(g9649,g2227,g2153);
  nor NOR_19551(g9664,g4878,g4871,g4864,g4836);
  nor NOR_19552(g9694,g1936,g1862);
  nor NOR_19553(g9700,g2361,g2287);
  nor NOR_19554(g9755,g2070,g1996);
  nor NOR_19555(g9762,g2495,g2421);
  nor NOR_19556(g9835,g2629,g2555);
  nor NOR_19557(g10123,g4294,g4297);
  nor NOR_19558(g10179,g2098,g1964,g1830,g1696);
  nor NOR_19559(g10205,g2657,g2523,g2389,g2255);
  nor NOR_19560(g10266,g5188,g5180);
  nor NOR_19561(g10281,g5535,g5527);
  nor NOR_19562(g10312,g5881,g5873);
  nor NOR_19563(g10318,g25,g22);
  nor NOR_19564(g10338,g5062,g5022);
  nor NOR_19565(g10341,g6227,g6219);
  nor NOR_19566(g10421,g6227,g9518);
  nor NOR_19567(g10488,g4616,g7133,g10336);
  nor NOR_19568(g10491,g6573,g9576);
  nor NOR_19569(g10510,g7183,g4593,g4584);
  nor NOR_19570(g10555,g7227,g4601,g4608);
  nor NOR_19571(g10615,g1636,g7308);
  nor NOR_19572(g10649,g1183,g8407);
  nor NOR_19573(g10666,g8462,g1171);
  nor NOR_19574(g10671,g1526,g8466);
  nor NOR_19575(g10695,g8462,g8407);
  nor NOR_19576(g10699,g8526,g1514);
  nor NOR_19577(g10709,g7499,g351);
  nor NOR_19578(g10715,g8526,g8466);
  nor NOR_19579(g10760,g1046,g7479);
  nor NOR_19580(g10793,g1389,g7503);
  nor NOR_19581(g10799,g347,g7541);
  nor NOR_19582(g10801,g1041,g7479);
  nor NOR_19583(g10803,g1384,g7503);
  nor NOR_19584(g10808,g8509,g7611);
  nor NOR_19585(g10819,g7479,g1041);
  nor NOR_19586(g10821,g7503,g1384);
  nor NOR_19587(g10831,g7690,g7827);
  nor NOR_19588(g10862,g7701,g7840);
  nor NOR_19589(g10884,g7650,g8451);
  nor NOR_19590(g10893,g1189,g7715,g7749);
  nor NOR_19591(g10899,g4064,g8451);
  nor NOR_19592(g10918,g1532,g7751,g7778);
  nor NOR_19593(g10922,g7650,g4057);
  nor NOR_19594(g11006,g7686,g7836);
  nor NOR_19595(g11012,g7693,g7846);
  nor NOR_19596(g11039,g9056,g9092);
  nor NOR_19597(g11107,g9095,g9177);
  nor NOR_19598(g11119,g9180,g9203);
  nor NOR_19599(g11148,g8052,g9197,g9174,g9050);
  nor NOR_19600(g11171,g8088,g9226,g9200,g9091);
  nor NOR_19601(g11184,g513,g9040);
  nor NOR_19602(g11185,g8038,g8183,g6804);
  nor NOR_19603(g11191,g4776,g4801,g9030);
  nor NOR_19604(g11194,g3288,g6875);
  nor NOR_19605(g11201,g4125,g7765);
  nor NOR_19606(g11203,g4966,g4991,g9064);
  nor NOR_19607(g11207,g3639,g6905);
  nor NOR_19608(g11213,g4776,g7892,g9030);
  nor NOR_19609(g11216,g7998,g8037);
  nor NOR_19610(g11217,g8531,g6875);
  nor NOR_19611(g11225,g3990,g6928);
  nor NOR_19612(g11231,g7928,g4801,g4793);
  nor NOR_19613(g11232,g4966,g7898,g9064);
  nor NOR_19614(g11238,g8584,g6905);
  nor NOR_19615(g11248,g7953,g4991,g4983);
  nor NOR_19616(g11252,g8620,g3057);
  nor NOR_19617(g11255,g8623,g6928);
  nor NOR_19618(g11261,g7928,g4801,g9030);
  nor NOR_19619(g11270,g8431,g8434);
  nor NOR_19620(g11273,g3061,g8620);
  nor NOR_19621(g11276,g8534,g8691);
  nor NOR_19622(g11280,g8647,g3408);
  nor NOR_19623(g11283,g7953,g4991,g9064);
  nor NOR_19624(g11303,g8497,g8500);
  nor NOR_19625(g11306,g3412,g8647);
  nor NOR_19626(g11309,g8587,g8728);
  nor NOR_19627(g11313,g8669,g3759);
  nor NOR_19628(g11345,g8477,g8479);
  nor NOR_19629(g11346,g7980,g7964);
  nor NOR_19630(g11357,g8558,g8561);
  nor NOR_19631(g11360,g3763,g8669);
  nor NOR_19632(g11363,g8626,g8751);
  nor NOR_19633(g11384,g8538,g8540);
  nor NOR_19634(g11385,g8021,g7985);
  nor NOR_19635(g11414,g8591,g8593);
  nor NOR_19636(g11415,g8080,g8026);
  nor NOR_19637(g11435,g8107,g3171);
  nor NOR_19638(g11448,g4191,g8790);
  nor NOR_19639(g11469,g650,g9903,g645);
  nor NOR_19640(g11473,g8107,g8059);
  nor NOR_19641(g11483,g8165,g3522);
  nor NOR_19642(g11493,g8964,g8967);
  nor NOR_19643(g11514,g10295,g3161,g3155);
  nor NOR_19644(g11527,g8165,g8114);
  nor NOR_19645(g11537,g8229,g3873);
  nor NOR_19646(g11563,g8059,g8011);
  nor NOR_19647(g11566,g3161,g7964);
  nor NOR_19648(g11571,g10323,g3512,g3506);
  nor NOR_19649(g11584,g8229,g8172);
  nor NOR_19650(g11607,g8848,g8993,g376);
  nor NOR_19651(g11610,g7980,g3155);
  nor NOR_19652(g11618,g8114,g8070);
  nor NOR_19653(g11621,g3512,g7985);
  nor NOR_19654(g11626,g7121,g3863,g3857);
  nor NOR_19655(g11653,g7980,g7964);
  nor NOR_19656(g11658,g8021,g3506);
  nor NOR_19657(g11666,g8172,g8125);
  nor NOR_19658(g11669,g3863,g8026);
  nor NOR_19659(g11692,g8021,g7985);
  nor NOR_19660(g11697,g8080,g3857);
  nor NOR_19661(g11715,g8080,g8026);
  nor NOR_19662(g11729,g3179,g8059);
  nor NOR_19663(g11747,g3530,g8114);
  nor NOR_19664(g11755,g4709,g8796);
  nor NOR_19665(g11763,g3881,g8172);
  nor NOR_19666(g11771,g8921,g4185);
  nor NOR_19667(g11773,g8883,g4785);
  nor NOR_19668(g11780,g4899,g8822);
  nor NOR_19669(g11797,g8883,g8796);
  nor NOR_19670(g11804,g8938,g4975);
  nor NOR_19671(g11834,g8938,g8822);
  nor NOR_19672(g11846,g7635,g7518,g7548);
  nor NOR_19673(g11862,g7134,g7150);
  nor NOR_19674(g11869,g7649,g7534,g7581);
  nor NOR_19675(g11885,g7153,g7167);
  nor NOR_19676(g11891,g812,g9166);
  nor NOR_19677(g11907,g7170,g7184);
  nor NOR_19678(g11913,g7197,g9166);
  nor NOR_19679(g11924,g7187,g7209);
  nor NOR_19680(g11932,g843,g9166);
  nor NOR_19681(g11935,g9485,g7267);
  nor NOR_19682(g11940,g2712,g10084);
  nor NOR_19683(g11945,g7212,g7228);
  nor NOR_19684(g11950,g9220,g9166);
  nor NOR_19685(g11954,g9538,g7314);
  nor NOR_19686(g11958,g9543,g7327);
  nor NOR_19687(g11972,g9591,g7361);
  nor NOR_19688(g11976,g9595,g7379);
  nor NOR_19689(g11995,g9645,g7410);
  nor NOR_19690(g11999,g9654,g7423);
  nor NOR_19691(g12002,g5297,g7004);
  nor NOR_19692(g12017,g9969,g9586);
  nor NOR_19693(g12025,g9705,g7461);
  nor NOR_19694(g12026,g9417,g9340);
  nor NOR_19695(g12029,g5644,g7028);
  nor NOR_19696(g12046,g10036,g9640);
  nor NOR_19697(g12050,g10038,g9649);
  nor NOR_19698(g12059,g9853,g7004);
  nor NOR_19699(g12067,g5990,g7051);
  nor NOR_19700(g12081,g10079,g9694);
  nor NOR_19701(g12085,g10082,g9700);
  nor NOR_19702(g12093,g9924,g7028);
  nor NOR_19703(g12101,g6336,g7074);
  nor NOR_19704(g12113,g1648,g8187);
  nor NOR_19705(g12117,g10113,g9755);
  nor NOR_19706(g12121,g10117,g9762);
  nor NOR_19707(g12123,g6856,g2748);
  nor NOR_19708(g12126,g9989,g5069);
  nor NOR_19709(g12129,g9992,g7051);
  nor NOR_19710(g12137,g6682,g7097);
  nor NOR_19711(g12146,g1783,g8241);
  nor NOR_19712(g12150,g2208,g8259);
  nor NOR_19713(g12154,g10155,g9835);
  nor NOR_19714(g12160,g9721,g9724);
  nor NOR_19715(g12163,g5073,g9989);
  nor NOR_19716(g12166,g9856,g10124);
  nor NOR_19717(g12170,g10047,g5413);
  nor NOR_19718(g12173,g10050,g7074);
  nor NOR_19719(g12189,g1917,g8302);
  nor NOR_19720(g12193,g2342,g8316);
  nor NOR_19721(g12198,g9797,g9800);
  nor NOR_19722(g12201,g5417,g10047);
  nor NOR_19723(g12204,g9927,g10160);
  nor NOR_19724(g12208,g10096,g5759);
  nor NOR_19725(g12211,g10099,g7097);
  nor NOR_19726(g12223,g2051,g8365);
  nor NOR_19727(g12226,g2476,g8373);
  nor NOR_19728(g12228,g10222,g10206,g10184,g10335);
  nor NOR_19729(g12234,g9776,g9778);
  nor NOR_19730(g12235,g9234,g9206);
  nor NOR_19731(g12246,g9880,g9883);
  nor NOR_19732(g12249,g5763,g10096);
  nor NOR_19733(g12252,g9995,g10185);
  nor NOR_19734(g12256,g10136,g6105);
  nor NOR_19735(g12288,g2610,g8418);
  nor NOR_19736(g12296,g9860,g9862);
  nor NOR_19737(g12297,g9269,g9239);
  nor NOR_19738(g12308,g9951,g9954);
  nor NOR_19739(g12311,g6109,g10136);
  nor NOR_19740(g12314,g10053,g10207);
  nor NOR_19741(g12318,g10172,g6451);
  nor NOR_19742(g12333,g1624,g8139);
  nor NOR_19743(g12346,g9931,g9933);
  nor NOR_19744(g12347,g9321,g9274);
  nor NOR_19745(g12358,g10019,g10022);
  nor NOR_19746(g12361,g6455,g10172);
  nor NOR_19747(g12364,g10102,g10224);
  nor NOR_19748(g12371,g1760,g8195);
  nor NOR_19749(g12374,g2185,g8205);
  nor NOR_19750(g12377,g6856,g2748,g9708);
  nor NOR_19751(g12405,g9374,g5180);
  nor NOR_19752(g12418,g9999,g10001);
  nor NOR_19753(g12419,g9402,g9326);
  nor NOR_19754(g12432,g1894,g8249);
  nor NOR_19755(g12435,g9012,g8956,g8904,g8863);
  nor NOR_19756(g12437,g2319,g8267);
  nor NOR_19757(g12443,g9374,g9300);
  nor NOR_19758(g12453,g9444,g5527);
  nor NOR_19759(g12466,g10057,g10059);
  nor NOR_19760(g12467,g9472,g9407);
  nor NOR_19761(g12479,g2028,g8310);
  nor NOR_19762(g12483,g2453,g8324);
  nor NOR_19763(g12486,g9055,g9013,g8957,g8905);
  nor NOR_19764(g12492,g7704,g5170,g5164);
  nor NOR_19765(g12505,g9444,g9381);
  nor NOR_19766(g12515,g9511,g5873);
  nor NOR_19767(g12540,g2587,g8381);
  nor NOR_19768(g12550,g9300,g9259);
  nor NOR_19769(g12553,g5170,g9206);
  nor NOR_19770(g12558,g7738,g5517,g5511);
  nor NOR_19771(g12571,g9511,g9451);
  nor NOR_19772(g12581,g9569,g6219);
  nor NOR_19773(g12591,g504,g9040);
  nor NOR_19774(g12593,g9234,g5164);
  nor NOR_19775(g12601,g9381,g9311);
  nor NOR_19776(g12604,g5517,g9239);
  nor NOR_19777(g12609,g7766,g5863,g5857);
  nor NOR_19778(g12622,g9569,g9518);
  nor NOR_19779(g12632,g9631,g6565);
  nor NOR_19780(g12645,g4467,g6961);
  nor NOR_19781(g12646,g9234,g9206);
  nor NOR_19782(g12651,g9269,g5511);
  nor NOR_19783(g12659,g9451,g9392);
  nor NOR_19784(g12662,g5863,g9274);
  nor NOR_19785(g12667,g7791,g6209,g6203);
  nor NOR_19786(g12680,g9631,g9576);
  nor NOR_19787(g12695,g9269,g9239);
  nor NOR_19788(g12700,g9321,g5857);
  nor NOR_19789(g12708,g9518,g9462);
  nor NOR_19790(g12711,g6209,g9326);
  nor NOR_19791(g12716,g7812,g6555,g6549);
  nor NOR_19792(g12729,g1657,g8139);
  nor NOR_19793(g12739,g9321,g9274);
  nor NOR_19794(g12744,g9402,g6203);
  nor NOR_19795(g12752,g9576,g9529);
  nor NOR_19796(g12755,g6555,g9407);
  nor NOR_19797(g12772,g5188,g9300);
  nor NOR_19798(g12780,g9402,g9326);
  nor NOR_19799(g12785,g9472,g6549);
  nor NOR_19800(g12798,g5535,g9381);
  nor NOR_19801(g12806,g9472,g9407);
  nor NOR_19802(g12821,g7132,g10223,g7149,g10261);
  nor NOR_19803(g12824,g5881,g9451);
  nor NOR_19804(g12846,g6837,g10430);
  nor NOR_19805(g12847,g6838,g10430);
  nor NOR_19806(g12848,g6839,g10430);
  nor NOR_19807(g12849,g6840,g10430);
  nor NOR_19808(g12850,g10430,g6845);
  nor NOR_19809(g12851,g6846,g10430);
  nor NOR_19810(g12852,g6847,g10430);
  nor NOR_19811(g12853,g6848,g10430);
  nor NOR_19812(g12854,g6849,g10430);
  nor NOR_19813(g12855,g10430,g6854);
  nor NOR_19814(g12856,g10430,g6855);
  nor NOR_19815(g12858,g10365,g10430);
  nor NOR_19816(g12970,g10555,g10510,g10488);
  nor NOR_19817(g12980,g7909,g10741);
  nor NOR_19818(g13004,g7933,g10741);
  nor NOR_19819(g13005,g7939,g10762);
  nor NOR_19820(g13013,g7957,g10762);
  nor NOR_19821(g13021,g7544,g10741);
  nor NOR_19822(g13031,g7301,g10741);
  nor NOR_19823(g13032,g7577,g10762);
  nor NOR_19824(g13044,g7349,g10762);
  nor NOR_19825(g13056,g7400,g10741);
  nor NOR_19826(g13076,g7443,g10741);
  nor NOR_19827(g13078,g7446,g10762);
  nor NOR_19828(g13094,g7487,g10762);
  nor NOR_19829(g13110,g7841,g10741);
  nor NOR_19830(g13114,g7528,g10741);
  nor NOR_19831(g13125,g7863,g10762);
  nor NOR_19832(g13129,g7553,g10762);
  nor NOR_19833(g13202,g8347,g10511);
  nor NOR_19834(g13325,g7841,g10741);
  nor NOR_19835(g13326,g10929,g10905);
  nor NOR_19836(g13335,g7851,g10741);
  nor NOR_19837(g13336,g11330,g11011);
  nor NOR_19838(g13341,g7863,g10762);
  nor NOR_19839(g13342,g10961,g10935);
  nor NOR_19840(g13377,g7873,g10762);
  nor NOR_19841(g13378,g11374,g11017);
  nor NOR_19842(g13480,g3017,g11858);
  nor NOR_19843(g13500,g8480,g12641);
  nor NOR_19844(g13501,g3368,g11881);
  nor NOR_19845(g13512,g9077,g12527);
  nor NOR_19846(g13517,g8541,g12692);
  nor NOR_19847(g13518,g3719,g11903);
  nor NOR_19848(g13539,g8594,g12735);
  nor NOR_19849(g13568,g8046,g12527);
  nor NOR_19850(g13603,g8009,g10721);
  nor NOR_19851(g13622,g278,g11166);
  nor NOR_19852(g13631,g8068,g10733);
  nor NOR_19853(g13661,g528,g11185);
  nor NOR_19854(g13670,g8123,g10756);
  nor NOR_19855(g13698,g528,g12527,g11185);
  nor NOR_19856(g13700,g3288,g11615);
  nor NOR_19857(g13730,g3639,g11663);
  nor NOR_19858(g13765,g8531,g11615);
  nor NOR_19859(g13772,g3990,g11702);
  nor NOR_19860(g13796,g9158,g12527);
  nor NOR_19861(g13799,g8584,g11663);
  nor NOR_19862(g13806,g11245,g4076);
  nor NOR_19863(g13824,g8623,g11702);
  nor NOR_19864(g13831,g11245,g7666);
  nor NOR_19865(g13852,g11320,g8347);
  nor NOR_19866(g13872,g8745,g11083);
  nor NOR_19867(g13883,g4709,g4785,g11155);
  nor NOR_19868(g13908,g4709,g8796,g11155);
  nor NOR_19869(g13910,g4899,g4975,g11173);
  nor NOR_19870(g13913,g8859,g11083);
  nor NOR_19871(g13919,g3347,g11276);
  nor NOR_19872(g13937,g8883,g4785,g11155);
  nor NOR_19873(g13939,g4899,g8822,g11173);
  nor NOR_19874(g13944,g10262,g12259);
  nor NOR_19875(g13946,g8651,g11083);
  nor NOR_19876(g13947,g8948,g11083);
  nor NOR_19877(g13954,g8663,g11276);
  nor NOR_19878(g13959,g3698,g11309);
  nor NOR_19879(g13970,g8883,g8796,g11155);
  nor NOR_19880(g13971,g8938,g4975,g11173);
  nor NOR_19881(g13989,g8697,g11309);
  nor NOR_19882(g13994,g4049,g11363);
  nor NOR_19883(g13996,g8938,g8822,g11173);
  nor NOR_19884(g14000,g8766,g12259);
  nor NOR_19885(g14001,g739,g11083);
  nor NOR_19886(g14002,g8681,g11083);
  nor NOR_19887(g14003,g9003,g11083);
  nor NOR_19888(g14027,g8734,g11363);
  nor NOR_19889(g14033,g8808,g12259);
  nor NOR_19890(g14036,g8725,g11083);
  nor NOR_19891(g14037,g8748,g11083);
  nor NOR_19892(g14064,g9214,g12259);
  nor NOR_19893(g14090,g8851,g12259);
  nor NOR_19894(g14091,g8854,g12259);
  nor NOR_19895(g14092,g8774,g11083);
  nor NOR_19896(g14093,g8833,g11083);
  nor NOR_19897(g14094,g8770,g11083);
  nor NOR_19898(g14121,g8891,g12259);
  nor NOR_19899(g14122,g8895,g12259);
  nor NOR_19900(g14124,g8830,g11083);
  nor NOR_19901(g14145,g8945,g12259);
  nor NOR_19902(g14163,g8997,g12259);
  nor NOR_19903(g14164,g9000,g12259);
  nor NOR_19904(g14165,g8951,g11083);
  nor NOR_19905(g14176,g9044,g12259);
  nor NOR_19906(g14178,g8899,g11083);
  nor NOR_19907(g14181,g9083,g12259);
  nor NOR_19908(g14188,g9162,g12259);
  nor NOR_19909(g14194,g5029,g10515);
  nor NOR_19910(g14211,g9779,g10823);
  nor NOR_19911(g14212,g5373,g10537);
  nor NOR_19912(g14227,g9863,g10838);
  nor NOR_19913(g14228,g5719,g10561);
  nor NOR_19914(g14247,g9934,g10869);
  nor NOR_19915(g14248,g6065,g10578);
  nor NOR_19916(g14253,g10032,g12259,g9217);
  nor NOR_19917(g14271,g10002,g10874);
  nor NOR_19918(g14272,g6411,g10598);
  nor NOR_19919(g14278,g562,g12259,g9217);
  nor NOR_19920(g14291,g9839,g12155);
  nor NOR_19921(g14306,g10060,g10887);
  nor NOR_19922(g14313,g12016,g9250);
  nor NOR_19923(g14320,g9257,g11111);
  nor NOR_19924(g14334,g12044,g9337);
  nor NOR_19925(g14335,g12045,g9283);
  nor NOR_19926(g14337,g12049,g9284);
  nor NOR_19927(g14339,g12289,g2735);
  nor NOR_19928(g14347,g9309,g11123);
  nor NOR_19929(g14360,g12078,g9484);
  nor NOR_19930(g14361,g12079,g9413);
  nor NOR_19931(g14362,g12080,g9338);
  nor NOR_19932(g14364,g12083,g9415);
  nor NOR_19933(g14365,g12084,g9339);
  nor NOR_19934(g14367,g9547,g12289);
  nor NOR_19935(g14382,g9390,g11139);
  nor NOR_19936(g14391,g12112,g9585);
  nor NOR_19937(g14392,g12114,g9537);
  nor NOR_19938(g14393,g12115,g9488);
  nor NOR_19939(g14394,g12116,g9414);
  nor NOR_19940(g14395,g12118,g9542);
  nor NOR_19941(g14396,g12119,g9489);
  nor NOR_19942(g14397,g12120,g9416);
  nor NOR_19943(g14399,g5297,g12598);
  nor NOR_19944(g14411,g9460,g11160);
  nor NOR_19945(g14413,g11914,g9638);
  nor NOR_19946(g14414,g12145,g9639);
  nor NOR_19947(g14415,g12147,g9590);
  nor NOR_19948(g14416,g12148,g9541);
  nor NOR_19949(g14417,g12149,g9648);
  nor NOR_19950(g14418,g12151,g9594);
  nor NOR_19951(g14419,g12152,g9546);
  nor NOR_19952(g14420,g12153,g9490);
  nor NOR_19953(g14425,g5644,g12656);
  nor NOR_19954(g14437,g9527,g11178);
  nor NOR_19955(g14444,g11936,g9692);
  nor NOR_19956(g14445,g12188,g9693);
  nor NOR_19957(g14446,g12190,g9644);
  nor NOR_19958(g14447,g11938,g9698);
  nor NOR_19959(g14448,g12192,g9699);
  nor NOR_19960(g14449,g12194,g9653);
  nor NOR_19961(g14450,g12195,g9598);
  nor NOR_19962(g14490,g9853,g12598);
  nor NOR_19963(g14497,g5990,g12705);
  nor NOR_19964(g14512,g11955,g9753);
  nor NOR_19965(g14513,g12222,g9754);
  nor NOR_19966(g14514,g11959,g9760);
  nor NOR_19967(g14515,g12225,g9761);
  nor NOR_19968(g14516,g12227,g9704);
  nor NOR_19969(g14522,g9924,g12656);
  nor NOR_19970(g14529,g6336,g12749);
  nor NOR_19971(g14538,g11973,g9828);
  nor NOR_19972(g14539,g11977,g9833);
  nor NOR_19973(g14540,g12287,g9834);
  nor NOR_19974(g14549,g9992,g12705);
  nor NOR_19975(g14556,g6682,g12790);
  nor NOR_19976(g14568,g12000,g9915);
  nor NOR_19977(g14575,g10050,g12749);
  nor NOR_19978(g14602,g10099,g12790);
  nor NOR_19979(g14611,g12333,g9749);
  nor NOR_19980(g14640,g12371,g9824);
  nor NOR_19981(g14642,g12374,g9829);
  nor NOR_19982(g14678,g12432,g9907);
  nor NOR_19983(g14679,g12437,g9911);
  nor NOR_19984(g14687,g5352,g12166);
  nor NOR_19985(g14707,g10143,g12259);
  nor NOR_19986(g14712,g12479,g9971);
  nor NOR_19987(g14713,g12483,g9974);
  nor NOR_19988(g14726,g10090,g12166);
  nor NOR_19989(g14731,g5698,g12204);
  nor NOR_19990(g14751,g10622,g10617,g10609,g10603);
  nor NOR_19991(g14752,g12540,g10040);
  nor NOR_19992(g14754,g12821,g2988);
  nor NOR_19993(g14767,g10130,g12204);
  nor NOR_19994(g14772,g6044,g12252);
  nor NOR_19995(g14792,g10653,g10623,g10618,g10611);
  nor NOR_19996(g14793,g2988,g12228);
  nor NOR_19997(g14816,g10166,g12252);
  nor NOR_19998(g14821,g6390,g12314);
  nor NOR_19999(g14867,g10191,g12314);
  nor NOR_20000(g14872,g6736,g12364);
  nor NOR_20001(g14911,g10213,g12364);
  nor NOR_20002(g14914,g12822,g12797);
  nor NOR_20003(g14988,g10816,g10812,g10805);
  nor NOR_20004(g15049,g13350,g6799);
  nor NOR_20005(g15050,g12834,g13350);
  nor NOR_20006(g15051,g6801,g13350);
  nor NOR_20007(g15052,g12835,g13350);
  nor NOR_20008(g15053,g12836,g13350);
  nor NOR_20009(g15054,g12837,g13350);
  nor NOR_20010(g15055,g6808,g13350);
  nor NOR_20011(g15056,g6809,g13350);
  nor NOR_20012(g15057,g6810,g13350);
  nor NOR_20013(g15058,g12838,g13350);
  nor NOR_20014(g15059,g12839,g13350);
  nor NOR_20015(g15060,g13350,g6814);
  nor NOR_20016(g15061,g6815,g13394);
  nor NOR_20017(g15062,g6817,g13394);
  nor NOR_20018(g15063,g6818,g13394);
  nor NOR_20019(g15064,g6820,g13394);
  nor NOR_20020(g15065,g13394,g12840);
  nor NOR_20021(g15066,g12841,g13394);
  nor NOR_20022(g15067,g12842,g13394);
  nor NOR_20023(g15068,g6826,g13416);
  nor NOR_20024(g15069,g6828,g13416);
  nor NOR_20025(g15070,g6829,g13416);
  nor NOR_20026(g15071,g6831,g13416);
  nor NOR_20027(g15072,g13416,g12843);
  nor NOR_20028(g15073,g12844,g13416);
  nor NOR_20029(g15074,g12845,g13416);
  nor NOR_20030(g15086,g13144,g12859);
  nor NOR_20031(g15087,g12860,g13144);
  nor NOR_20032(g15088,g13144,g6874);
  nor NOR_20033(g15089,g13144,g12861);
  nor NOR_20034(g15090,g13144,g12862);
  nor NOR_20035(g15091,g13177,g12863);
  nor NOR_20036(g15092,g12864,g13177);
  nor NOR_20037(g15093,g13177,g6904);
  nor NOR_20038(g15094,g13177,g12865);
  nor NOR_20039(g15095,g13177,g12866);
  nor NOR_20040(g15096,g13191,g12867);
  nor NOR_20041(g15097,g12868,g13191);
  nor NOR_20042(g15098,g13191,g6927);
  nor NOR_20043(g15099,g13191,g12869);
  nor NOR_20044(g15100,g13191,g12870);
  nor NOR_20045(g15101,g12871,g14591);
  nor NOR_20046(g15102,g14591,g6954);
  nor NOR_20047(g15106,g12872,g10430);
  nor NOR_20048(g15120,g12873,g13605);
  nor NOR_20049(g15121,g12874,g13605);
  nor NOR_20050(g15122,g6959,g13605);
  nor NOR_20051(g15123,g6975,g13605);
  nor NOR_20052(g15126,g12878,g13605);
  nor NOR_20053(g15127,g12879,g13605);
  nor NOR_20054(g15128,g13638,g12880);
  nor NOR_20055(g15129,g6984,g13638);
  nor NOR_20056(g15130,g13638,g6985);
  nor NOR_20057(g15131,g12881,g13638);
  nor NOR_20058(g15132,g12882,g13638);
  nor NOR_20059(g15133,g12883,g13638);
  nor NOR_20060(g15134,g13638,g12884);
  nor NOR_20061(g15135,g6990,g13638);
  nor NOR_20062(g15136,g13680,g12885);
  nor NOR_20063(g15137,g6992,g13680);
  nor NOR_20064(g15138,g13680,g6993);
  nor NOR_20065(g15139,g12886,g13680);
  nor NOR_20066(g15140,g12887,g13680);
  nor NOR_20067(g15141,g12888,g13680);
  nor NOR_20068(g15142,g13680,g12889);
  nor NOR_20069(g15143,g6998,g13680);
  nor NOR_20070(g15144,g13716,g12890);
  nor NOR_20071(g15145,g12891,g13716);
  nor NOR_20072(g15146,g13716,g7003);
  nor NOR_20073(g15147,g13716,g12892);
  nor NOR_20074(g15148,g13716,g12893);
  nor NOR_20075(g15149,g13745,g12894);
  nor NOR_20076(g15150,g12895,g13745);
  nor NOR_20077(g15151,g13745,g7027);
  nor NOR_20078(g15152,g13745,g12896);
  nor NOR_20079(g15153,g13745,g12897);
  nor NOR_20080(g15154,g13782,g12898);
  nor NOR_20081(g15155,g12899,g13782);
  nor NOR_20082(g15156,g13782,g7050);
  nor NOR_20083(g15157,g13782,g12900);
  nor NOR_20084(g15158,g13782,g12901);
  nor NOR_20085(g15159,g13809,g12902);
  nor NOR_20086(g15160,g12903,g13809);
  nor NOR_20087(g15161,g13809,g7073);
  nor NOR_20088(g15162,g13809,g12904);
  nor NOR_20089(g15163,g13809,g12905);
  nor NOR_20090(g15164,g13835,g12906);
  nor NOR_20091(g15165,g12907,g13835);
  nor NOR_20092(g15166,g13835,g7096);
  nor NOR_20093(g15167,g13835,g12908);
  nor NOR_20094(g15168,g13835,g12909);
  nor NOR_20095(g15170,g7118,g14279);
  nor NOR_20096(g15372,g817,g14279);
  nor NOR_20097(g15508,g10320,g14279);
  nor NOR_20098(g15570,g822,g14279);
  nor NOR_20099(g15578,g7216,g14279);
  nor NOR_20100(g15585,g11862,g14194);
  nor NOR_20101(g15594,g10614,g13026,g7285);
  nor NOR_20102(g15608,g11885,g14212);
  nor NOR_20103(g15628,g11907,g14228);
  nor NOR_20104(g15647,g11924,g14248);
  nor NOR_20105(g15669,g11945,g14272);
  nor NOR_20106(g15718,g13858,g11330);
  nor NOR_20107(g15724,g13858,g11374);
  nor NOR_20108(g15754,g341,g7440,g13385);
  nor NOR_20109(g15825,g7666,g13217);
  nor NOR_20110(g15992,g10929,g13846);
  nor NOR_20111(g16024,g14216,g11890);
  nor NOR_20112(g16027,g10929,g13260);
  nor NOR_20113(g16044,g10961,g13861);
  nor NOR_20114(g16066,g10929,g13307);
  nor NOR_20115(g16072,g10961,g13273);
  nor NOR_20116(g16090,g10961,g13315);
  nor NOR_20117(g16183,g9223,g13545);
  nor NOR_20118(g16198,g9247,g13574);
  nor NOR_20119(g16201,g13462,g4704);
  nor NOR_20120(g16209,g13478,g4749);
  nor NOR_20121(g16210,g13479,g4894);
  nor NOR_20122(g16215,g1211,g13545);
  nor NOR_20123(g16219,g13498,g4760);
  nor NOR_20124(g16220,g13499,g4939);
  nor NOR_20125(g16226,g8052,g13545);
  nor NOR_20126(g16227,g1554,g13574);
  nor NOR_20127(g16231,g13515,g4771);
  nor NOR_20128(g16232,g13516,g4950);
  nor NOR_20129(g16237,g8088,g13574);
  nor NOR_20130(g16242,g13529,g4961);
  nor NOR_20131(g16246,g13551,g11169);
  nor NOR_20132(g16268,g7913,g13121);
  nor NOR_20133(g16272,g13580,g11189);
  nor NOR_20134(g16287,g13622,g11144);
  nor NOR_20135(g16288,g13794,g417);
  nor NOR_20136(g16292,g7943,g13134);
  nor NOR_20137(g16313,g8005,g13600);
  nor NOR_20138(g16424,g8064,g13628);
  nor NOR_20139(g16476,g8119,g13667);
  nor NOR_20140(g16479,g14719,g12490);
  nor NOR_20141(g16488,g13697,g13656);
  nor NOR_20142(g16581,g13756,g8086);
  nor NOR_20143(g16646,g13437,g11020,g11372);
  nor NOR_20144(g17148,g827,g14279);
  nor NOR_20145(g17174,g9194,g14279);
  nor NOR_20146(g17175,g1216,g13545);
  nor NOR_20147(g17180,g1559,g13574);
  nor NOR_20148(g17190,g723,g14279);
  nor NOR_20149(g17194,g11039,g13480);
  nor NOR_20150(g17198,g9282,g14279);
  nor NOR_20151(g17213,g11107,g13501);
  nor NOR_20152(g17239,g11119,g13518);
  nor NOR_20153(g17284,g9253,g14317);
  nor NOR_20154(g17309,g9305,g14344);
  nor NOR_20155(g17393,g9386,g14379);
  nor NOR_20156(g17420,g9456,g14408);
  nor NOR_20157(g17482,g9523,g14434);
  nor NOR_20158(g17515,g13221,g10828);
  nor NOR_20159(g17619,g10179,g12955);
  nor NOR_20160(g17625,g14541,g12123);
  nor NOR_20161(g17657,g14751,g12955);
  nor NOR_20162(g17663,g10205,g12983);
  nor NOR_20163(g17694,g12435,g12955);
  nor NOR_20164(g17700,g14792,g12983);
  nor NOR_20165(g17727,g12486,g12983);
  nor NOR_20166(g17954,g832,g14279);
  nor NOR_20167(g19063,g7909,g15674);
  nor NOR_20168(g19070,g16957,g11720);
  nor NOR_20169(g19140,g7939,g15695);
  nor NOR_20170(g19209,g12971,g15614,g11320);
  nor NOR_20171(g19268,g15979,g962);
  nor NOR_20172(g19338,g16031,g1306);
  nor NOR_20173(g19388,g17181,g14256);
  nor NOR_20174(g19400,g17139,g14206);
  nor NOR_20175(g19401,g17193,g14296);
  nor NOR_20176(g19402,g15979,g13133);
  nor NOR_20177(g19413,g17151,g14221);
  nor NOR_20178(g19422,g16031,g13141);
  nor NOR_20179(g19430,g17150,g14220);
  nor NOR_20180(g19436,g17176,g14233);
  nor NOR_20181(g19444,g17192,g14295);
  nor NOR_20182(g19453,g17199,g14316);
  nor NOR_20183(g19778,g16268,g1061);
  nor NOR_20184(g19793,g16292,g1404);
  nor NOR_20185(g19853,g15746,g1052);
  nor NOR_20186(g19873,g15755,g1395);
  nor NOR_20187(g19880,g16201,g13634);
  nor NOR_20188(g19887,g3025,g16275);
  nor NOR_20189(g19890,g16987,g8058);
  nor NOR_20190(g19906,g16209,g13672);
  nor NOR_20191(g19907,g16210,g13676);
  nor NOR_20192(g19919,g16987,g11205);
  nor NOR_20193(g19932,g3376,g16296);
  nor NOR_20194(g19935,g17062,g8113);
  nor NOR_20195(g19951,g16219,g13709);
  nor NOR_20196(g19953,g16220,g13712);
  nor NOR_20197(g19968,g17062,g11223);
  nor NOR_20198(g19981,g3727,g16316);
  nor NOR_20199(g19984,g17096,g8171);
  nor NOR_20200(g19997,g16231,g13739);
  nor NOR_20201(g19999,g16232,g13742);
  nor NOR_20202(g20000,g13661,g16264);
  nor NOR_20203(g20014,g17096,g11244);
  nor NOR_20204(g20027,g16242,g13779);
  nor NOR_20205(g20149,g17091,g14185);
  nor NOR_20206(g20183,g17152,g14222);
  nor NOR_20207(g20234,g17140,g14207);
  nor NOR_20208(g20390,g17182,g14257);
  nor NOR_20209(g20717,g5037,g17217);
  nor NOR_20210(g20720,g17847,g9299);
  nor NOR_20211(g20841,g17847,g12027);
  nor NOR_20212(g20854,g5381,g17243);
  nor NOR_20213(g20857,g17929,g9380);
  nor NOR_20214(g20982,g17929,g12065);
  nor NOR_20215(g20995,g5727,g17287);
  nor NOR_20216(g20998,g18065,g9450);
  nor NOR_20217(g21062,g9547,g17297);
  nor NOR_20218(g21127,g18065,g12099);
  nor NOR_20219(g21140,g6073,g17312);
  nor NOR_20220(g21143,g15348,g9517);
  nor NOR_20221(g21193,g15348,g12135);
  nor NOR_20222(g21206,g6419,g17396);
  nor NOR_20223(g21209,g15483,g9575);
  nor NOR_20224(g21250,g9417,g9340,g17494);
  nor NOR_20225(g21256,g15483,g12179);
  nor NOR_20226(g21277,g9417,g9340,g17467);
  nor NOR_20227(g21284,g16646,g9690);
  nor NOR_20228(g21389,g10143,g17748,g12259);
  nor NOR_20229(g21652,g17619,g17663);
  nor NOR_20230(g21655,g17657,g17700);
  nor NOR_20231(g21658,g17694,g17727);
  nor NOR_20232(g22190,g2827,g18949);
  nor NOR_20233(g22357,g1024,g19699);
  nor NOR_20234(g22399,g1367,g19720);
  nor NOR_20235(g22400,g19345,g15718);
  nor NOR_20236(g22405,g18957,g20136,g20114);
  nor NOR_20237(g22448,g1018,g19699);
  nor NOR_20238(g22450,g19345,g15724);
  nor NOR_20239(g22488,g19699,g1002);
  nor NOR_20240(g22491,g1361,g19720);
  nor NOR_20241(g22513,g1002,g19699);
  nor NOR_20242(g22514,g19699,g1018);
  nor NOR_20243(g22517,g19720,g1345);
  nor NOR_20244(g22521,g1036,g19699);
  nor NOR_20245(g22522,g19699,g1024);
  nor NOR_20246(g22523,g1345,g19720);
  nor NOR_20247(g22524,g19720,g1361);
  nor NOR_20248(g22535,g19699,g1030);
  nor NOR_20249(g22536,g1379,g19720);
  nor NOR_20250(g22537,g19720,g1367);
  nor NOR_20251(g22539,g1030,g19699);
  nor NOR_20252(g22540,g19720,g1373);
  nor NOR_20253(g22545,g1373,g19720);
  nor NOR_20254(g22654,g7733,g19506);
  nor NOR_20255(g22929,g19773,g12970);
  nor NOR_20256(g22983,g979,g16268,g19853);
  nor NOR_20257(g22993,g1322,g16292,g19873);
  nor NOR_20258(g23024,g7936,g19407);
  nor NOR_20259(g23042,g16581,g19462,g10685);
  nor NOR_20260(g23051,g7960,g19427);
  nor NOR_20261(g23052,g8334,g19916);
  nor NOR_20262(g23063,g16313,g19887);
  nor NOR_20263(g23079,g8390,g19965);
  nor NOR_20264(g23108,g16424,g19932);
  nor NOR_20265(g23124,g8443,g20011);
  nor NOR_20266(g23135,g16476,g19981);
  nor NOR_20267(g23204,g10685,g19462,g16488);
  nor NOR_20268(g23208,g20035,g16324);
  nor NOR_20269(g23560,g9607,g20838);
  nor NOR_20270(g23586,g17284,g20717);
  nor NOR_20271(g23602,g9672,g20979);
  nor NOR_20272(g23626,g17309,g20854);
  nor NOR_20273(g23642,g9733,g21124);
  nor NOR_20274(g23662,g17393,g20995);
  nor NOR_20275(g23678,g9809,g21190);
  nor NOR_20276(g23686,g2767,g21066);
  nor NOR_20277(g23695,g17420,g21140);
  nor NOR_20278(g23711,g9892,g21253);
  nor NOR_20279(g23729,g17482,g21206);
  nor NOR_20280(g23763,g2795,g21276);
  nor NOR_20281(g23835,g2791,g21303);
  nor NOR_20282(g23871,g2811,g21348);
  nor NOR_20283(g23883,g2779,g21067);
  nor NOR_20284(g23918,g2799,g21382);
  nor NOR_20285(g23955,g2823,g18890);
  nor NOR_20286(g23956,g18957,g18918,g20136,g20114);
  nor NOR_20287(g24018,I23162,I23163);
  nor NOR_20288(g24145,g19402,g19422);
  nor NOR_20289(g24148,g19268,g19338);
  nor NOR_20290(g24383,g22409,g22360);
  nor NOR_20291(g24391,g22190,g14645);
  nor NOR_20292(g24439,g7400,g22312);
  nor NOR_20293(g24453,g7446,g22325);
  nor NOR_20294(g24494,g23513,g23532);
  nor NOR_20295(g24497,g23533,g23553);
  nor NOR_20296(g24508,g23577,g23618);
  nor NOR_20297(g24514,g23619,g23657);
  nor NOR_20298(g24575,g23498,g23514);
  nor NOR_20299(g24619,g23554,g23581);
  nor NOR_20300(g24631,g20516,g20436,g20219,g22957);
  nor NOR_20301(g24701,g979,g23024,g19778);
  nor NOR_20302(g24720,g1322,g23051,g19793);
  nor NOR_20303(g24751,g3034,g23105);
  nor NOR_20304(g24766,g3385,g23132);
  nor NOR_20305(g24779,g3736,g23167);
  nor NOR_20306(g24875,g8725,g23850,g11083);
  nor NOR_20307(g24953,g10262,g23978,g12259);
  nor NOR_20308(g24959,g8858,g23324);
  nor NOR_20309(g24976,g671,g23324);
  nor NOR_20310(g24990,g8898,g23324);
  nor NOR_20311(g25004,g676,g23324);
  nor NOR_20312(g25005,g6811,g23324);
  nor NOR_20313(g25022,g714,g23324);
  nor NOR_20314(g25141,g22228,g10334);
  nor NOR_20315(g25144,g5046,g23623);
  nor NOR_20316(g25160,g5390,g23659);
  nor NOR_20317(g25175,g5736,g23692);
  nor NOR_20318(g25189,g6082,g23726);
  nor NOR_20319(g25203,g6428,g23756);
  nor NOR_20320(g25247,g23763,g14645);
  nor NOR_20321(g25317,g9766,g23782);
  nor NOR_20322(g25321,g23835,g14645);
  nor NOR_20323(g25407,g23871,g14645);
  nor NOR_20324(g25446,g23686,g14645);
  nor NOR_20325(g25447,g23883,g14645);
  nor NOR_20326(g25501,g23918,g14645);
  nor NOR_20327(g25504,g22550,g7222);
  nor NOR_20328(g25521,g23955,g14645);
  nor NOR_20329(g25540,g22409,g22360);
  nor NOR_20330(g25769,g25453,g25414);
  nor NOR_20331(g25770,g25417,g25377);
  nor NOR_20332(g25776,g7166,g24380,g24369);
  nor NOR_20333(g25777,g25482,g25456);
  nor NOR_20334(g25778,g25459,g25420);
  nor NOR_20335(g25784,g25507,g25485);
  nor NOR_20336(g25785,g25488,g25462);
  nor NOR_20337(g25800,g25518,g25510);
  nor NOR_20338(g25851,g4311,g24380,g24369);
  nor NOR_20339(g25887,g24984,g11706);
  nor NOR_20340(g25932,g7680,g24528);
  nor NOR_20341(g25944,g7716,g24591);
  nor NOR_20342(g25947,g1199,g24591);
  nor NOR_20343(g25948,g7752,g24609);
  nor NOR_20344(g25950,g1070,g24591);
  nor NOR_20345(g25952,g1542,g24609);
  nor NOR_20346(g25954,g7750,g24591);
  nor NOR_20347(g25956,g1413,g24609);
  nor NOR_20348(g25958,g7779,g24609);
  nor NOR_20349(g26098,g9073,g24732);
  nor NOR_20350(g26162,g23052,g24751);
  nor NOR_20351(g26183,g23079,g24766);
  nor NOR_20352(g26209,g23124,g24779);
  nor NOR_20353(g26212,g23837,g25408);
  nor NOR_20354(g26247,g7995,g24732);
  nor NOR_20355(g26256,g23873,g25479);
  nor NOR_20356(g26267,g8033,g24732);
  nor NOR_20357(g26268,g283,g24825);
  nor NOR_20358(g26296,g8287,g24732);
  nor NOR_20359(g26297,g8519,g24825);
  nor NOR_20360(g26298,g8297,g24825);
  nor NOR_20361(g26309,g8575,g24825);
  nor NOR_20362(g26314,g24808,g24802);
  nor NOR_20363(g26330,g8631,g24825);
  nor NOR_20364(g26338,g8458,g24825);
  nor NOR_20365(g26346,g8522,g24825);
  nor NOR_20366(g26515,g24843,g24822);
  nor NOR_20367(g26545,g24881,g24855);
  nor NOR_20368(g26546,g24858,g24846);
  nor NOR_20369(g26573,g24897,g24884);
  nor NOR_20370(g26574,g24887,g24861);
  nor NOR_20371(g26598,g8990,g13756,g24732);
  nor NOR_20372(g26603,g24908,g24900);
  nor NOR_20373(g26609,g146,g24732);
  nor NOR_20374(g26625,g23560,g25144);
  nor NOR_20375(g26628,g8990,g24732);
  nor NOR_20376(g26645,g23602,g25160);
  nor NOR_20377(g26649,g9037,g24732);
  nor NOR_20378(g26667,g23642,g25175);
  nor NOR_20379(g26686,g23678,g25189);
  nor NOR_20380(g26715,g23711,g25203);
  nor NOR_20381(g26865,g25328,g25290);
  nor NOR_20382(g26872,g25411,g25371);
  nor NOR_20383(g26873,g25374,g25331);
  nor NOR_20384(g26976,g5016,g25791);
  nor NOR_20385(g26993,g5360,g25805);
  nor NOR_20386(g27007,g5706,g25821);
  nor NOR_20387(g27010,g6052,g25839);
  nor NOR_20388(g27012,g6398,g25856);
  nor NOR_20389(g27027,g26398,g26484);
  nor NOR_20390(g27046,g7544,g25888);
  nor NOR_20391(g27059,g7577,g25895);
  nor NOR_20392(g27063,g26485,g26516);
  nor NOR_20393(g27093,g26712,g26749);
  nor NOR_20394(g27102,g26750,g26779);
  nor NOR_20395(g27337,g8334,g26616);
  nor NOR_20396(g27338,g9291,g26616);
  nor NOR_20397(g27343,g8005,g26616);
  nor NOR_20398(g27344,g8390,g26636);
  nor NOR_20399(g27345,g9360,g26636);
  nor NOR_20400(g27352,g7975,g26616);
  nor NOR_20401(g27353,g8097,g26616);
  nor NOR_20402(g27354,g8064,g26636);
  nor NOR_20403(g27355,g8443,g26657);
  nor NOR_20404(g27356,g9429,g26657);
  nor NOR_20405(g27364,g8426,g26616);
  nor NOR_20406(g27366,g8016,g26636);
  nor NOR_20407(g27367,g8155,g26636);
  nor NOR_20408(g27368,g8119,g26657);
  nor NOR_20409(g27379,g8492,g26636);
  nor NOR_20410(g27381,g8075,g26657);
  nor NOR_20411(g27382,g8219,g26657);
  nor NOR_20412(g27400,g8553,g26657);
  nor NOR_20413(g27479,g9056,g26616);
  nor NOR_20414(g27499,g9095,g26636);
  nor NOR_20415(g27511,g22137,g26866,g20277);
  nor NOR_20416(g27516,g9180,g26657);
  nor NOR_20417(g27528,g8770,g26352,g11083);
  nor NOR_20418(g27629,g8891,g26382,g12259);
  nor NOR_20419(g27647,g3004,g26616);
  nor NOR_20420(g27652,g3355,g26636);
  nor NOR_20421(g27659,g3706,g26657);
  nor NOR_20422(g27703,g9607,g25791);
  nor NOR_20423(g27704,g7239,g25791);
  nor NOR_20424(g27717,g9492,g26745);
  nor NOR_20425(g27720,g9253,g25791);
  nor NOR_20426(g27721,g9672,g25805);
  nor NOR_20427(g27722,g7247,g25805);
  nor NOR_20428(g27731,g9229,g25791);
  nor NOR_20429(g27732,g9364,g25791);
  nor NOR_20430(g27733,g9305,g25805);
  nor NOR_20431(g27734,g9733,g25821);
  nor NOR_20432(g27735,g7262,g25821);
  nor NOR_20433(g27766,g9716,g25791);
  nor NOR_20434(g27768,g9264,g25805);
  nor NOR_20435(g27769,g9434,g25805);
  nor NOR_20436(g27770,g9386,g25821);
  nor NOR_20437(g27771,g9809,g25839);
  nor NOR_20438(g27772,g7297,g25839);
  nor NOR_20439(g27823,g9792,g25805);
  nor NOR_20440(g27825,g9316,g25821);
  nor NOR_20441(g27826,g9501,g25821);
  nor NOR_20442(g27827,g9456,g25839);
  nor NOR_20443(g27828,g9892,g25856);
  nor NOR_20444(g27829,g7345,g25856);
  nor NOR_20445(g27875,g9875,g25821);
  nor NOR_20446(g27877,g9397,g25839);
  nor NOR_20447(g27878,g9559,g25839);
  nor NOR_20448(g27879,g9523,g25856);
  nor NOR_20449(g27924,g9946,g25839);
  nor NOR_20450(g27926,g9467,g25856);
  nor NOR_20451(g27927,g9621,g25856);
  nor NOR_20452(g27954,g10014,g25856);
  nor NOR_20453(g27960,g7134,g25791);
  nor NOR_20454(g27966,g7153,g25805);
  nor NOR_20455(g27969,g7170,g25821);
  nor NOR_20456(g27973,g7187,g25839);
  nor NOR_20457(g27982,g7212,g25856);
  nor NOR_20458(g28031,g21209,I26522,I26523);
  nor NOR_20459(g28106,g7812,g26994);
  nor NOR_20460(g28149,g27598,g27612);
  nor NOR_20461(g28340,g27439,g26339);
  nor NOR_20462(g28353,g9073,g27654,g24732);
  nor NOR_20463(g28414,g27467,g26347);
  nor NOR_20464(g28425,g27493,g26351);
  nor NOR_20465(g28444,g8575,g27463,g24825);
  nor NOR_20466(g28452,g3161,g27602);
  nor NOR_20467(g28457,g7980,g27602);
  nor NOR_20468(g28462,g3512,g27617);
  nor NOR_20469(g28468,g3155,g10295,g27602);
  nor NOR_20470(g28469,g3171,g27602);
  nor NOR_20471(g28470,g8021,g27617);
  nor NOR_20472(g28475,g3863,g27635);
  nor NOR_20473(g28476,g27627,g26547);
  nor NOR_20474(g28480,g8059,g27602);
  nor NOR_20475(g28481,g3506,g10323,g27617);
  nor NOR_20476(g28482,g3522,g27617);
  nor NOR_20477(g28483,g8080,g27635);
  nor NOR_20478(g28491,g8114,g27617);
  nor NOR_20479(g28492,g3857,g7121,g27635);
  nor NOR_20480(g28493,g3873,g27635);
  nor NOR_20481(g28496,g3179,g27602);
  nor NOR_20482(g28498,g8172,g27635);
  nor NOR_20483(g28509,g8107,g27602);
  nor NOR_20484(g28510,g3530,g27617);
  nor NOR_20485(g28514,g8165,g27617);
  nor NOR_20486(g28515,g3881,g27635);
  nor NOR_20487(g28519,g8011,g27602,g10295);
  nor NOR_20488(g28520,g8229,g27635);
  nor NOR_20489(g28521,g27649,g26604);
  nor NOR_20490(g28529,g8070,g27617,g10323);
  nor NOR_20491(g28540,g8125,g27635,g7121);
  nor NOR_20492(g28552,g10295,g27602);
  nor NOR_20493(g28568,g10323,g27617);
  nor NOR_20494(g28584,g7121,g27635);
  nor NOR_20495(g28803,g27730,g22763);
  nor NOR_20496(g28953,g5170,g27999);
  nor NOR_20497(g28981,g9234,g27999);
  nor NOR_20498(g28986,g5517,g28010);
  nor NOR_20499(g29005,g5164,g7704,g27999);
  nor NOR_20500(g29006,g5180,g27999);
  nor NOR_20501(g29007,g9269,g28010);
  nor NOR_20502(g29012,g5863,g28020);
  nor NOR_20503(g29032,g9300,g27999);
  nor NOR_20504(g29033,g5511,g7738,g28010);
  nor NOR_20505(g29034,g5527,g28010);
  nor NOR_20506(g29035,g9321,g28020);
  nor NOR_20507(g29040,g6209,g26977);
  nor NOR_20508(g29069,g9381,g28010);
  nor NOR_20509(g29070,g5857,g7766,g28020);
  nor NOR_20510(g29071,g5873,g28020);
  nor NOR_20511(g29072,g9402,g26977);
  nor NOR_20512(g29077,g6555,g26994);
  nor NOR_20513(g29104,g5188,g27999);
  nor NOR_20514(g29106,g9451,g28020);
  nor NOR_20515(g29107,g6203,g7791,g26977);
  nor NOR_20516(g29108,g6219,g26977);
  nor NOR_20517(g29109,g9472,g26994);
  nor NOR_20518(g29141,g9374,g27999);
  nor NOR_20519(g29142,g5535,g28010);
  nor NOR_20520(g29144,g9518,g26977);
  nor NOR_20521(g29145,g6549,g7812,g26994);
  nor NOR_20522(g29146,g6565,g26994);
  nor NOR_20523(g29164,g9444,g28010);
  nor NOR_20524(g29165,g5881,g28020);
  nor NOR_20525(g29167,g9576,g26994);
  nor NOR_20526(g29173,g9259,g27999,g7704);
  nor NOR_20527(g29174,g9511,g28020);
  nor NOR_20528(g29175,g6227,g26977);
  nor NOR_20529(g29179,g9311,g28010,g7738);
  nor NOR_20530(g29180,g9569,g26977);
  nor NOR_20531(g29181,g6573,g26994);
  nor NOR_20532(g29183,g9392,g28020,g7766);
  nor NOR_20533(g29184,g9631,g26994);
  nor NOR_20534(g29187,g7704,g27999);
  nor NOR_20535(g29189,g9462,g26977,g7791);
  nor NOR_20536(g29191,g7738,g28010);
  nor NOR_20537(g29193,g9529,g26994,g7812);
  nor NOR_20538(g29198,g7766,g28020);
  nor NOR_20539(g29200,g7791,g26977);
  nor NOR_20540(g29359,g7528,g28167);
  nor NOR_20541(g29361,g7553,g28174);
  nor NOR_20542(g29370,g28585,g28599);
  nor NOR_20543(g29497,g22763,g28241);
  nor NOR_20544(g29503,g22763,g28250);
  nor NOR_20545(g29675,g28380,g8236,g8354);
  nor NOR_20546(g29705,g28399,g8284,g8404);
  nor NOR_20547(g29873,g6875,g28458);
  nor NOR_20548(g29886,g3288,g28458);
  nor NOR_20549(g29889,g6905,g28471);
  nor NOR_20550(g29898,g6895,g28458);
  nor NOR_20551(g29900,g3639,g28471);
  nor NOR_20552(g29903,g6928,g28484);
  nor NOR_20553(g29908,g6918,g28471);
  nor NOR_20554(g29910,g3990,g28484);
  nor NOR_20555(g29915,g6941,g28484);
  nor NOR_20556(g29916,g8681,g28504,g11083);
  nor NOR_20557(g29933,g8808,g28500,g12259);
  nor NOR_20558(g30106,g28739,g7268);
  nor NOR_20559(g30117,g28739,g7252);
  nor NOR_20560(g30119,g28761,g7315);
  nor NOR_20561(g30123,g28768,g7328);
  nor NOR_20562(g30129,g28739,g14537);
  nor NOR_20563(g30130,g28761,g7275);
  nor NOR_20564(g30132,g28789,g7362);
  nor NOR_20565(g30134,g28768,g7280);
  nor NOR_20566(g30136,g28799,g7380);
  nor NOR_20567(g30143,g28761,g14566);
  nor NOR_20568(g30144,g28789,g7322);
  nor NOR_20569(g30146,g28833,g7411);
  nor NOR_20570(g30147,g28768,g14567);
  nor NOR_20571(g30148,g28799,g7335);
  nor NOR_20572(g30150,g28846,g7424);
  nor NOR_20573(g30156,g28789,g14587);
  nor NOR_20574(g30157,g28833,g7369);
  nor NOR_20575(g30159,g28799,g14589);
  nor NOR_20576(g30160,g28846,g7387);
  nor NOR_20577(g30162,g28880,g7462);
  nor NOR_20578(g30169,g28833,g14613);
  nor NOR_20579(g30170,g28846,g14615);
  nor NOR_20580(g30171,g28880,g7431);
  nor NOR_20581(g30183,g28880,g14644);
  nor NOR_20582(g30240,g7004,g28982);
  nor NOR_20583(g30249,g5297,g28982);
  nor NOR_20584(g30252,g7028,g29008);
  nor NOR_20585(g30260,g7018,g28982);
  nor NOR_20586(g30262,g5644,g29008);
  nor NOR_20587(g30265,g7051,g29036);
  nor NOR_20588(g30271,g7041,g29008);
  nor NOR_20589(g30273,g5990,g29036);
  nor NOR_20590(g30276,g7074,g29073);
  nor NOR_20591(g30280,g7064,g29036);
  nor NOR_20592(g30282,g6336,g29073);
  nor NOR_20593(g30285,g7097,g29110);
  nor NOR_20594(g30288,g7087,g29073);
  nor NOR_20595(g30290,g6682,g29110);
  nor NOR_20596(g30294,g7110,g29110);
  nor NOR_20597(g30601,g16279,g29718);
  nor NOR_20598(g30613,g4507,g29365);
  nor NOR_20599(g30922,g16662,g29810);
  nor NOR_20600(g30929,g29803,g29835);
  nor NOR_20601(g30934,g29836,g29850);
  nor NOR_20602(g31008,g30004,g30026);
  nor NOR_20603(g31068,g4801,g29540);
  nor NOR_20604(g31116,g7892,g29540);
  nor NOR_20605(g31117,g4991,g29556);
  nor NOR_20606(g31119,g7898,g29556);
  nor NOR_20607(g31121,g4776,g29540);
  nor NOR_20608(g31126,g7928,g29540);
  nor NOR_20609(g31127,g4966,g29556);
  nor NOR_20610(g31133,g7953,g29556);
  nor NOR_20611(g31134,g8033,g29679,g24732);
  nor NOR_20612(g31233,g8522,g29778,g24825);
  nor NOR_20613(g31294,g11326,g29660);
  nor NOR_20614(g31318,g4785,g29697);
  nor NOR_20615(g31372,g8796,g29697);
  nor NOR_20616(g31373,g4975,g29725);
  nor NOR_20617(g31469,g8822,g29725);
  nor NOR_20618(g31476,g4709,g29697);
  nor NOR_20619(g31482,g8883,g29697);
  nor NOR_20620(g31483,g4899,g29725);
  nor NOR_20621(g31491,g8938,g29725);
  nor NOR_20622(g31498,g9030,g29540);
  nor NOR_20623(g31506,g4793,g29540);
  nor NOR_20624(g31507,g9064,g29556);
  nor NOR_20625(g31515,g4983,g29556);
  nor NOR_20626(g31935,g30583,g4349);
  nor NOR_20627(g31942,g8977,g30583);
  nor NOR_20628(g31965,g30583,g4358);
  nor NOR_20629(g31970,g9024,g30583);
  nor NOR_20630(g32017,g31504,g23475);
  nor NOR_20631(g32212,g8859,g31262,g11083);
  nor NOR_20632(g32296,g9044,g31509,g12259);
  nor NOR_20633(g32424,g8721,g31294);
  nor NOR_20634(g32455,g31566,I29985,I29986);
  nor NOR_20635(g32520,g31554,I30054,I30055);
  nor NOR_20636(g32585,g31542,I30123,I30124);
  nor NOR_20637(g32650,g31579,I30192,I30193);
  nor NOR_20638(g32715,g31327,I30261,I30262);
  nor NOR_20639(g32780,g31327,I30330,I30331);
  nor NOR_20640(g32845,g30673,I30399,I30400);
  nor NOR_20641(g32910,g31327,I30468,I30469);
  nor NOR_20642(g33075,g31997,g7163);
  nor NOR_20643(g33084,g31978,g7655);
  nor NOR_20644(g33085,g31978,g4311);
  nor NOR_20645(g33088,g31997,g7224);
  nor NOR_20646(g33089,g31978,g4322);
  nor NOR_20647(g33090,g31997,g4593);
  nor NOR_20648(g33092,g31978,g4332);
  nor NOR_20649(g33093,g31997,g4601);
  nor NOR_20650(g33094,g31950,g4639);
  nor NOR_20651(g33095,g31997,g7236);
  nor NOR_20652(g33096,g31997,g4608);
  nor NOR_20653(g33097,g31950,g4628);
  nor NOR_20654(g33098,g31997,g4616);
  nor NOR_20655(g33100,g32172,g31188);
  nor NOR_20656(g33103,g32176,g31212);
  nor NOR_20657(g33107,g32180,g31223);
  nor NOR_20658(g33108,g32183,g31228);
  nor NOR_20659(g33109,g31997,g4584);
  nor NOR_20660(g33112,g31240,g32194);
  nor NOR_20661(g33117,g31261,g32205);
  nor NOR_20662(g33125,g8606,g32057);
  nor NOR_20663(g33128,g4653,g32057);
  nor NOR_20664(g33129,g8630,g32072);
  nor NOR_20665(g33130,g32265,g31497);
  nor NOR_20666(g33131,g4659,g32057);
  nor NOR_20667(g33132,g4843,g32072);
  nor NOR_20668(g33133,g32278,g31503);
  nor NOR_20669(g33134,g7686,g32057);
  nor NOR_20670(g33135,g32090,g8350);
  nor NOR_20671(g33137,g4849,g32072);
  nor NOR_20672(g33138,g32287,g31514);
  nor NOR_20673(g33139,g8650,g32057);
  nor NOR_20674(g33140,g7693,g32072);
  nor NOR_20675(g33141,g32099,g8400);
  nor NOR_20676(g33143,g32293,g31518);
  nor NOR_20677(g33144,g4664,g32057);
  nor NOR_20678(g33145,g8677,g32072);
  nor NOR_20679(g33146,g4669,g32057);
  nor NOR_20680(g33147,g32090,g7788);
  nor NOR_20681(g33148,g4854,g32072);
  nor NOR_20682(g33160,g8672,g32057);
  nor NOR_20683(g33161,g32090,g7806);
  nor NOR_20684(g33162,g4859,g32072);
  nor NOR_20685(g33163,g32099,g7809);
  nor NOR_20686(g33174,g8714,g32072);
  nor NOR_20687(g33175,g32099,g7828);
  nor NOR_20688(g33419,g31978,g7627);
  nor NOR_20689(g33427,g10278,g31950);
  nor NOR_20690(g33432,g31997,g6978);
  nor NOR_20691(g33437,g31997,g10275);
  nor NOR_20692(g33438,g31950,g4621);
  nor NOR_20693(g33439,g31950,g4633);
  nor NOR_20694(g33447,g31978,g7643);
  nor NOR_20695(g33448,g7785,g31950);
  nor NOR_20696(g33449,g10311,g31950);
  nor NOR_20697(g33823,g8774,g33306,g11083);
  nor NOR_20698(g33851,g8854,g33299,g12259);
  nor NOR_20699(g34067,g33859,g11772);
  nor NOR_20700(g34354,g9003,g34162,g11083);
  nor NOR_20701(g34359,g9162,g34174,g12259);
  nor NOR_20702(g34496,g34370,g27648);
  nor NOR_20703(g34703,g8899,g34545,g11083);
  nor NOR_20704(g34737,g34706,g30003);
  nor NOR_20705(g34912,g34883,g20277,g20242,g21370);

endmodule