/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:00:16 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module AD42M1N ( CO, ICO, S, A, B, C, D, ICI );
   input A, B, C, D, ICI;
   output CO, ICO, S;
      AD42M1N_UDP5(CO, A, B, C, D, ICI);
      AD42M1N_UDP6(ICO, A, B, C);
      AD42M1N_UDP7(S, A, B, C, D, ICI);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO
    if (B===1'b0 && C===1'b0 && D===1'b0 && ICI===1'b1) 
        (A => CO) = (1.0, 1.0);
    if (B===1'b0 && C===1'b0 && D===1'b1 && ICI===1'b0) 
        (A => CO) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b1) 
        (A => CO) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b0) 
        (A => CO) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b1) 
        (A => CO) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b0) 
        (A => CO) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1 && D===1'b0 && ICI===1'b1) 
        (A => CO) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1 && D===1'b1 && ICI===1'b0) 
        (A => CO) = (1.0, 1.0);
    ifnone
        ( posedge A => ( CO +: A ) ) = (1.0, 1.0);
        ( negedge A => ( CO +: A ) ) = (1.0, 1.0);

    // arc A --> ICO
    if (B===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b0) 
        (A => ICO) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b1) 
        (A => ICO) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b0) 
        (A => ICO) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b1) 
        (A => ICO) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b0) 
        (A => ICO) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b1) 
        (A => ICO) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b0) 
        (A => ICO) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b1) 
        (A => ICO) = (1.0, 1.0);
    ifnone
        (A => ICO) = (1.0, 1.0);

    // arc A --> S
    if (B===1'b0 && C===1'b0 && D===1'b0 && ICI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && C===1'b0 && D===1'b0 && ICI===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && C===1'b0 && D===1'b1 && ICI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && C===1'b0 && D===1'b1 && ICI===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1 && D===1'b0 && ICI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1 && D===1'b0 && ICI===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1 && D===1'b1 && ICI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1 && D===1'b1 && ICI===1'b1) 
        (A => S) = (1.0, 1.0);
    ifnone
        ( posedge A => ( S +: A ) ) = (1.0, 1.0);
        ( negedge A => ( S +: A ) ) = (1.0, 1.0);

    // arc B --> CO
    if (A===1'b0 && C===1'b0 && D===1'b0 && ICI===1'b1) 
        (B => CO) = (1.0, 1.0);
    if (A===1'b0 && C===1'b0 && D===1'b1 && ICI===1'b0) 
        (B => CO) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b1) 
        (B => CO) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b0) 
        (B => CO) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b1) 
        (B => CO) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b0) 
        (B => CO) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1 && D===1'b0 && ICI===1'b1) 
        (B => CO) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1 && D===1'b1 && ICI===1'b0) 
        (B => CO) = (1.0, 1.0);
    ifnone
        ( posedge B => ( CO +: B ) ) = (1.0, 1.0);
        ( negedge B => ( CO +: B ) ) = (1.0, 1.0);

    // arc B --> ICO
    if (A===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b0) 
        (B => ICO) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b1) 
        (B => ICO) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b0) 
        (B => ICO) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b1) 
        (B => ICO) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b0) 
        (B => ICO) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b1) 
        (B => ICO) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b0) 
        (B => ICO) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b1) 
        (B => ICO) = (1.0, 1.0);
    ifnone
        (B => ICO) = (1.0, 1.0);

    // arc B --> S
    if (A===1'b0 && C===1'b0 && D===1'b0 && ICI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && C===1'b0 && D===1'b0 && ICI===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && C===1'b0 && D===1'b1 && ICI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && C===1'b0 && D===1'b1 && ICI===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1 && D===1'b0 && ICI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1 && D===1'b0 && ICI===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1 && D===1'b1 && ICI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1 && D===1'b1 && ICI===1'b1) 
        (B => S) = (1.0, 1.0);
    ifnone
        ( posedge B => ( S +: B ) ) = (1.0, 1.0);
        ( negedge B => ( S +: B ) ) = (1.0, 1.0);

    // arc C --> CO
    if (A===1'b0 && B===1'b0 && D===1'b0 && ICI===1'b1) 
        (C => CO) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && D===1'b1 && ICI===1'b0) 
        (C => CO) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && D===1'b0 && ICI===1'b1) 
        (C => CO) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && D===1'b1 && ICI===1'b0) 
        (C => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && D===1'b0 && ICI===1'b1) 
        (C => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && D===1'b1 && ICI===1'b0) 
        (C => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && D===1'b0 && ICI===1'b1) 
        (C => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && D===1'b1 && ICI===1'b0) 
        (C => CO) = (1.0, 1.0);
    ifnone
        ( posedge C => ( CO +: C ) ) = (1.0, 1.0);
        ( negedge C => ( CO +: C ) ) = (1.0, 1.0);

    // arc C --> ICO
    if (A===1'b0 && B===1'b1 && D===1'b0 && ICI===1'b0) 
        (C => ICO) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && D===1'b0 && ICI===1'b1) 
        (C => ICO) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && D===1'b1 && ICI===1'b0) 
        (C => ICO) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && D===1'b1 && ICI===1'b1) 
        (C => ICO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && D===1'b0 && ICI===1'b0) 
        (C => ICO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && D===1'b0 && ICI===1'b1) 
        (C => ICO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && D===1'b1 && ICI===1'b0) 
        (C => ICO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && D===1'b1 && ICI===1'b1) 
        (C => ICO) = (1.0, 1.0);
    ifnone
        (C => ICO) = (1.0, 1.0);

    // arc C --> S
    if (A===1'b0 && B===1'b0 && D===1'b0 && ICI===1'b0) 
        (C => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && D===1'b0 && ICI===1'b1) 
        (C => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && D===1'b1 && ICI===1'b0) 
        (C => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && D===1'b1 && ICI===1'b1) 
        (C => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && D===1'b0 && ICI===1'b0) 
        (C => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && D===1'b0 && ICI===1'b1) 
        (C => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && D===1'b1 && ICI===1'b0) 
        (C => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && D===1'b1 && ICI===1'b1) 
        (C => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && D===1'b0 && ICI===1'b0) 
        (C => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && D===1'b0 && ICI===1'b1) 
        (C => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && D===1'b1 && ICI===1'b0) 
        (C => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && D===1'b1 && ICI===1'b1) 
        (C => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && D===1'b0 && ICI===1'b0) 
        (C => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && D===1'b0 && ICI===1'b1) 
        (C => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && D===1'b1 && ICI===1'b0) 
        (C => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && D===1'b1 && ICI===1'b1) 
        (C => S) = (1.0, 1.0);
    ifnone
        ( posedge C => ( S +: C ) ) = (1.0, 1.0);
        ( negedge C => ( S +: C ) ) = (1.0, 1.0);

    // arc D --> CO
    if (A===1'b0 && B===1'b0 && C===1'b0 && ICI===1'b1) 
        (D => CO) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && ICI===1'b0) 
        (D => CO) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && ICI===1'b0) 
        (D => CO) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && ICI===1'b1) 
        (D => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && ICI===1'b0) 
        (D => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && ICI===1'b1) 
        (D => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && ICI===1'b1) 
        (D => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && ICI===1'b0) 
        (D => CO) = (1.0, 1.0);
    ifnone
        (D => CO) = (1.0, 1.0);

    // arc D --> S
    if (A===1'b0 && B===1'b0 && C===1'b0 && ICI===1'b0) 
        (D => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b0 && ICI===1'b1) 
        (D => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && ICI===1'b0) 
        (D => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && ICI===1'b1) 
        (D => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && ICI===1'b0) 
        (D => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && ICI===1'b1) 
        (D => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && ICI===1'b0) 
        (D => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && ICI===1'b1) 
        (D => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && ICI===1'b0) 
        (D => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && ICI===1'b1) 
        (D => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && ICI===1'b0) 
        (D => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && ICI===1'b1) 
        (D => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && ICI===1'b0) 
        (D => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && ICI===1'b1) 
        (D => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && ICI===1'b0) 
        (D => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && ICI===1'b1) 
        (D => S) = (1.0, 1.0);
    ifnone
        ( posedge D => ( S +: D ) ) = (1.0, 1.0);
        ( negedge D => ( S +: D ) ) = (1.0, 1.0);

    // arc ICI --> CO
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1) 
        (ICI => CO) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0) 
        (ICI => CO) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0) 
        (ICI => CO) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1) 
        (ICI => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0) 
        (ICI => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1) 
        (ICI => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1) 
        (ICI => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0) 
        (ICI => CO) = (1.0, 1.0);
    ifnone
        (ICI => CO) = (1.0, 1.0);

    // arc ICI --> S
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b0) 
        (ICI => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1) 
        (ICI => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0) 
        (ICI => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1) 
        (ICI => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0) 
        (ICI => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1) 
        (ICI => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0) 
        (ICI => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1) 
        (ICI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0) 
        (ICI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1) 
        (ICI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0) 
        (ICI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1) 
        (ICI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0) 
        (ICI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1) 
        (ICI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0) 
        (ICI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b1) 
        (ICI => S) = (1.0, 1.0);
    ifnone
        ( posedge ICI => ( S +: ICI ) ) = (1.0, 1.0);
        ( negedge ICI => ( S +: ICI ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AD42M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:00:31 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module AD42M2N ( CO, ICO, S, A, B, C, D, ICI );
   input A, B, C, D, ICI;
   output CO, ICO, S;
      AD42M1N_UDP5(CO, A, B, C, D, ICI);
      AD42M1N_UDP6(ICO, A, B, C);
      AD42M1N_UDP7(S, A, B, C, D, ICI);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO
    if (B===1'b0 && C===1'b0 && D===1'b0 && ICI===1'b1) 
        (A => CO) = (1.0, 1.0);
    if (B===1'b0 && C===1'b0 && D===1'b1 && ICI===1'b0) 
        (A => CO) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b1) 
        (A => CO) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b0) 
        (A => CO) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b1) 
        (A => CO) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b0) 
        (A => CO) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1 && D===1'b0 && ICI===1'b1) 
        (A => CO) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1 && D===1'b1 && ICI===1'b0) 
        (A => CO) = (1.0, 1.0);
    ifnone
        ( posedge A => ( CO +: A ) ) = (1.0, 1.0);
        ( negedge A => ( CO +: A ) ) = (1.0, 1.0);

    // arc A --> ICO
    if (B===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b0) 
        (A => ICO) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b1) 
        (A => ICO) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b0) 
        (A => ICO) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b1) 
        (A => ICO) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b0) 
        (A => ICO) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b1) 
        (A => ICO) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b0) 
        (A => ICO) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b1) 
        (A => ICO) = (1.0, 1.0);
    ifnone
        (A => ICO) = (1.0, 1.0);

    // arc A --> S
    if (B===1'b0 && C===1'b0 && D===1'b0 && ICI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && C===1'b0 && D===1'b0 && ICI===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && C===1'b0 && D===1'b1 && ICI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && C===1'b0 && D===1'b1 && ICI===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1 && D===1'b0 && ICI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1 && D===1'b0 && ICI===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1 && D===1'b1 && ICI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1 && D===1'b1 && ICI===1'b1) 
        (A => S) = (1.0, 1.0);
    ifnone
        ( posedge A => ( S +: A ) ) = (1.0, 1.0);
        ( negedge A => ( S +: A ) ) = (1.0, 1.0);

    // arc B --> CO
    if (A===1'b0 && C===1'b0 && D===1'b0 && ICI===1'b1) 
        (B => CO) = (1.0, 1.0);
    if (A===1'b0 && C===1'b0 && D===1'b1 && ICI===1'b0) 
        (B => CO) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b1) 
        (B => CO) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b0) 
        (B => CO) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b1) 
        (B => CO) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b0) 
        (B => CO) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1 && D===1'b0 && ICI===1'b1) 
        (B => CO) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1 && D===1'b1 && ICI===1'b0) 
        (B => CO) = (1.0, 1.0);
    ifnone
        ( posedge B => ( CO +: B ) ) = (1.0, 1.0);
        ( negedge B => ( CO +: B ) ) = (1.0, 1.0);

    // arc B --> ICO
    if (A===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b0) 
        (B => ICO) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b1) 
        (B => ICO) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b0) 
        (B => ICO) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b1) 
        (B => ICO) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b0) 
        (B => ICO) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b1) 
        (B => ICO) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b0) 
        (B => ICO) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b1) 
        (B => ICO) = (1.0, 1.0);
    ifnone
        (B => ICO) = (1.0, 1.0);

    // arc B --> S
    if (A===1'b0 && C===1'b0 && D===1'b0 && ICI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && C===1'b0 && D===1'b0 && ICI===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && C===1'b0 && D===1'b1 && ICI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && C===1'b0 && D===1'b1 && ICI===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1 && D===1'b0 && ICI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1 && D===1'b0 && ICI===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1 && D===1'b1 && ICI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1 && D===1'b1 && ICI===1'b1) 
        (B => S) = (1.0, 1.0);
    ifnone
        ( posedge B => ( S +: B ) ) = (1.0, 1.0);
        ( negedge B => ( S +: B ) ) = (1.0, 1.0);

    // arc C --> CO
    if (A===1'b0 && B===1'b0 && D===1'b0 && ICI===1'b1) 
        (C => CO) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && D===1'b1 && ICI===1'b0) 
        (C => CO) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && D===1'b0 && ICI===1'b1) 
        (C => CO) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && D===1'b1 && ICI===1'b0) 
        (C => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && D===1'b0 && ICI===1'b1) 
        (C => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && D===1'b1 && ICI===1'b0) 
        (C => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && D===1'b0 && ICI===1'b1) 
        (C => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && D===1'b1 && ICI===1'b0) 
        (C => CO) = (1.0, 1.0);
    ifnone
        ( posedge C => ( CO +: C ) ) = (1.0, 1.0);
        ( negedge C => ( CO +: C ) ) = (1.0, 1.0);

    // arc C --> ICO
    if (A===1'b0 && B===1'b1 && D===1'b0 && ICI===1'b0) 
        (C => ICO) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && D===1'b0 && ICI===1'b1) 
        (C => ICO) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && D===1'b1 && ICI===1'b0) 
        (C => ICO) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && D===1'b1 && ICI===1'b1) 
        (C => ICO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && D===1'b0 && ICI===1'b0) 
        (C => ICO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && D===1'b0 && ICI===1'b1) 
        (C => ICO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && D===1'b1 && ICI===1'b0) 
        (C => ICO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && D===1'b1 && ICI===1'b1) 
        (C => ICO) = (1.0, 1.0);
    ifnone
        (C => ICO) = (1.0, 1.0);

    // arc C --> S
    if (A===1'b0 && B===1'b0 && D===1'b0 && ICI===1'b0) 
        (C => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && D===1'b0 && ICI===1'b1) 
        (C => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && D===1'b1 && ICI===1'b0) 
        (C => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && D===1'b1 && ICI===1'b1) 
        (C => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && D===1'b0 && ICI===1'b0) 
        (C => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && D===1'b0 && ICI===1'b1) 
        (C => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && D===1'b1 && ICI===1'b0) 
        (C => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && D===1'b1 && ICI===1'b1) 
        (C => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && D===1'b0 && ICI===1'b0) 
        (C => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && D===1'b0 && ICI===1'b1) 
        (C => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && D===1'b1 && ICI===1'b0) 
        (C => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && D===1'b1 && ICI===1'b1) 
        (C => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && D===1'b0 && ICI===1'b0) 
        (C => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && D===1'b0 && ICI===1'b1) 
        (C => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && D===1'b1 && ICI===1'b0) 
        (C => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && D===1'b1 && ICI===1'b1) 
        (C => S) = (1.0, 1.0);
    ifnone
        ( posedge C => ( S +: C ) ) = (1.0, 1.0);
        ( negedge C => ( S +: C ) ) = (1.0, 1.0);

    // arc D --> CO
    if (A===1'b0 && B===1'b0 && C===1'b0 && ICI===1'b1) 
        (D => CO) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && ICI===1'b0) 
        (D => CO) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && ICI===1'b0) 
        (D => CO) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && ICI===1'b1) 
        (D => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && ICI===1'b0) 
        (D => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && ICI===1'b1) 
        (D => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && ICI===1'b1) 
        (D => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && ICI===1'b0) 
        (D => CO) = (1.0, 1.0);
    ifnone
        (D => CO) = (1.0, 1.0);

    // arc D --> S
    if (A===1'b0 && B===1'b0 && C===1'b0 && ICI===1'b0) 
        (D => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b0 && ICI===1'b1) 
        (D => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && ICI===1'b0) 
        (D => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && ICI===1'b1) 
        (D => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && ICI===1'b0) 
        (D => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && ICI===1'b1) 
        (D => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && ICI===1'b0) 
        (D => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && ICI===1'b1) 
        (D => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && ICI===1'b0) 
        (D => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && ICI===1'b1) 
        (D => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && ICI===1'b0) 
        (D => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && ICI===1'b1) 
        (D => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && ICI===1'b0) 
        (D => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && ICI===1'b1) 
        (D => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && ICI===1'b0) 
        (D => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && ICI===1'b1) 
        (D => S) = (1.0, 1.0);
    ifnone
        ( posedge D => ( S +: D ) ) = (1.0, 1.0);
        ( negedge D => ( S +: D ) ) = (1.0, 1.0);

    // arc ICI --> CO
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1) 
        (ICI => CO) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0) 
        (ICI => CO) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0) 
        (ICI => CO) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1) 
        (ICI => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0) 
        (ICI => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1) 
        (ICI => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1) 
        (ICI => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0) 
        (ICI => CO) = (1.0, 1.0);
    ifnone
        (ICI => CO) = (1.0, 1.0);

    // arc ICI --> S
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b0) 
        (ICI => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1) 
        (ICI => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0) 
        (ICI => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1) 
        (ICI => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0) 
        (ICI => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1) 
        (ICI => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0) 
        (ICI => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1) 
        (ICI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0) 
        (ICI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1) 
        (ICI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0) 
        (ICI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1) 
        (ICI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0) 
        (ICI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1) 
        (ICI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0) 
        (ICI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b1) 
        (ICI => S) = (1.0, 1.0);
    ifnone
        ( posedge ICI => ( S +: ICI ) ) = (1.0, 1.0);
        ( negedge ICI => ( S +: ICI ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AD42M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:01:15 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module AD42M4N ( CO, ICO, S, A, B, C, D, ICI );
   input A, B, C, D, ICI;
   output CO, ICO, S;
      AD42M1N_UDP5(CO, A, B, C, D, ICI);
      AD42M1N_UDP6(ICO, A, B, C);
      AD42M1N_UDP7(S, A, B, C, D, ICI);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO
    if (B===1'b0 && C===1'b0 && D===1'b0 && ICI===1'b1) 
        (A => CO) = (1.0, 1.0);
    if (B===1'b0 && C===1'b0 && D===1'b1 && ICI===1'b0) 
        (A => CO) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b1) 
        (A => CO) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b0) 
        (A => CO) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b1) 
        (A => CO) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b0) 
        (A => CO) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1 && D===1'b0 && ICI===1'b1) 
        (A => CO) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1 && D===1'b1 && ICI===1'b0) 
        (A => CO) = (1.0, 1.0);
    ifnone
        ( posedge A => ( CO +: A ) ) = (1.0, 1.0);
        ( negedge A => ( CO +: A ) ) = (1.0, 1.0);

    // arc A --> ICO
    if (B===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b0) 
        (A => ICO) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b1) 
        (A => ICO) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b0) 
        (A => ICO) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b1) 
        (A => ICO) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b0) 
        (A => ICO) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b1) 
        (A => ICO) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b0) 
        (A => ICO) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b1) 
        (A => ICO) = (1.0, 1.0);
    ifnone
        (A => ICO) = (1.0, 1.0);

    // arc A --> S
    if (B===1'b0 && C===1'b0 && D===1'b0 && ICI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && C===1'b0 && D===1'b0 && ICI===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && C===1'b0 && D===1'b1 && ICI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && C===1'b0 && D===1'b1 && ICI===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1 && D===1'b0 && ICI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1 && D===1'b0 && ICI===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1 && D===1'b1 && ICI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1 && D===1'b1 && ICI===1'b1) 
        (A => S) = (1.0, 1.0);
    ifnone
        ( posedge A => ( S +: A ) ) = (1.0, 1.0);
        ( negedge A => ( S +: A ) ) = (1.0, 1.0);

    // arc B --> CO
    if (A===1'b0 && C===1'b0 && D===1'b0 && ICI===1'b1) 
        (B => CO) = (1.0, 1.0);
    if (A===1'b0 && C===1'b0 && D===1'b1 && ICI===1'b0) 
        (B => CO) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b1) 
        (B => CO) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b0) 
        (B => CO) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b1) 
        (B => CO) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b0) 
        (B => CO) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1 && D===1'b0 && ICI===1'b1) 
        (B => CO) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1 && D===1'b1 && ICI===1'b0) 
        (B => CO) = (1.0, 1.0);
    ifnone
        ( posedge B => ( CO +: B ) ) = (1.0, 1.0);
        ( negedge B => ( CO +: B ) ) = (1.0, 1.0);

    // arc B --> ICO
    if (A===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b0) 
        (B => ICO) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b1) 
        (B => ICO) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b0) 
        (B => ICO) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b1) 
        (B => ICO) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b0) 
        (B => ICO) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b1) 
        (B => ICO) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b0) 
        (B => ICO) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b1) 
        (B => ICO) = (1.0, 1.0);
    ifnone
        (B => ICO) = (1.0, 1.0);

    // arc B --> S
    if (A===1'b0 && C===1'b0 && D===1'b0 && ICI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && C===1'b0 && D===1'b0 && ICI===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && C===1'b0 && D===1'b1 && ICI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && C===1'b0 && D===1'b1 && ICI===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1 && D===1'b0 && ICI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1 && D===1'b0 && ICI===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1 && D===1'b1 && ICI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1 && D===1'b1 && ICI===1'b1) 
        (B => S) = (1.0, 1.0);
    ifnone
        ( posedge B => ( S +: B ) ) = (1.0, 1.0);
        ( negedge B => ( S +: B ) ) = (1.0, 1.0);

    // arc C --> CO
    if (A===1'b0 && B===1'b0 && D===1'b0 && ICI===1'b1) 
        (C => CO) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && D===1'b1 && ICI===1'b0) 
        (C => CO) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && D===1'b0 && ICI===1'b1) 
        (C => CO) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && D===1'b1 && ICI===1'b0) 
        (C => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && D===1'b0 && ICI===1'b1) 
        (C => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && D===1'b1 && ICI===1'b0) 
        (C => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && D===1'b0 && ICI===1'b1) 
        (C => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && D===1'b1 && ICI===1'b0) 
        (C => CO) = (1.0, 1.0);
    ifnone
        ( posedge C => ( CO +: C ) ) = (1.0, 1.0);
        ( negedge C => ( CO +: C ) ) = (1.0, 1.0);

    // arc C --> ICO
    if (A===1'b0 && B===1'b1 && D===1'b0 && ICI===1'b0) 
        (C => ICO) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && D===1'b0 && ICI===1'b1) 
        (C => ICO) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && D===1'b1 && ICI===1'b0) 
        (C => ICO) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && D===1'b1 && ICI===1'b1) 
        (C => ICO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && D===1'b0 && ICI===1'b0) 
        (C => ICO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && D===1'b0 && ICI===1'b1) 
        (C => ICO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && D===1'b1 && ICI===1'b0) 
        (C => ICO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && D===1'b1 && ICI===1'b1) 
        (C => ICO) = (1.0, 1.0);
    ifnone
        (C => ICO) = (1.0, 1.0);

    // arc C --> S
    if (A===1'b0 && B===1'b0 && D===1'b0 && ICI===1'b0) 
        (C => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && D===1'b0 && ICI===1'b1) 
        (C => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && D===1'b1 && ICI===1'b0) 
        (C => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && D===1'b1 && ICI===1'b1) 
        (C => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && D===1'b0 && ICI===1'b0) 
        (C => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && D===1'b0 && ICI===1'b1) 
        (C => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && D===1'b1 && ICI===1'b0) 
        (C => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && D===1'b1 && ICI===1'b1) 
        (C => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && D===1'b0 && ICI===1'b0) 
        (C => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && D===1'b0 && ICI===1'b1) 
        (C => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && D===1'b1 && ICI===1'b0) 
        (C => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && D===1'b1 && ICI===1'b1) 
        (C => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && D===1'b0 && ICI===1'b0) 
        (C => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && D===1'b0 && ICI===1'b1) 
        (C => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && D===1'b1 && ICI===1'b0) 
        (C => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && D===1'b1 && ICI===1'b1) 
        (C => S) = (1.0, 1.0);
    ifnone
        ( posedge C => ( S +: C ) ) = (1.0, 1.0);
        ( negedge C => ( S +: C ) ) = (1.0, 1.0);

    // arc D --> CO
    if (A===1'b0 && B===1'b0 && C===1'b0 && ICI===1'b1) 
        (D => CO) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && ICI===1'b0) 
        (D => CO) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && ICI===1'b0) 
        (D => CO) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && ICI===1'b1) 
        (D => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && ICI===1'b0) 
        (D => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && ICI===1'b1) 
        (D => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && ICI===1'b1) 
        (D => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && ICI===1'b0) 
        (D => CO) = (1.0, 1.0);
    ifnone
        (D => CO) = (1.0, 1.0);

    // arc D --> S
    if (A===1'b0 && B===1'b0 && C===1'b0 && ICI===1'b0) 
        (D => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b0 && ICI===1'b1) 
        (D => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && ICI===1'b0) 
        (D => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && ICI===1'b1) 
        (D => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && ICI===1'b0) 
        (D => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && ICI===1'b1) 
        (D => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && ICI===1'b0) 
        (D => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && ICI===1'b1) 
        (D => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && ICI===1'b0) 
        (D => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && ICI===1'b1) 
        (D => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && ICI===1'b0) 
        (D => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && ICI===1'b1) 
        (D => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && ICI===1'b0) 
        (D => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && ICI===1'b1) 
        (D => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && ICI===1'b0) 
        (D => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && ICI===1'b1) 
        (D => S) = (1.0, 1.0);
    ifnone
        ( posedge D => ( S +: D ) ) = (1.0, 1.0);
        ( negedge D => ( S +: D ) ) = (1.0, 1.0);

    // arc ICI --> CO
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1) 
        (ICI => CO) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0) 
        (ICI => CO) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0) 
        (ICI => CO) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1) 
        (ICI => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0) 
        (ICI => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1) 
        (ICI => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1) 
        (ICI => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0) 
        (ICI => CO) = (1.0, 1.0);
    ifnone
        (ICI => CO) = (1.0, 1.0);

    // arc ICI --> S
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b0) 
        (ICI => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1) 
        (ICI => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0) 
        (ICI => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1) 
        (ICI => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0) 
        (ICI => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1) 
        (ICI => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0) 
        (ICI => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1) 
        (ICI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0) 
        (ICI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1) 
        (ICI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0) 
        (ICI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1) 
        (ICI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0) 
        (ICI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1) 
        (ICI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0) 
        (ICI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b1) 
        (ICI => S) = (1.0, 1.0);
    ifnone
        ( posedge ICI => ( S +: ICI ) ) = (1.0, 1.0);
        ( negedge ICI => ( S +: ICI ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AD42M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:05:09 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module ADCSCM2N ( CO0, CO1, A, B, NCI0, NCI1 );
   input A, B, NCI0, NCI1;
   output CO0, CO1;
      ADCSCM2N_UDP4(CO0, A, B, NCI0);
      ADCSCM2N_UDP5(CO1, A, B, NCI1);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO0
    if (B===1'b0 && NCI0===1'b0 && NCI1===1'b0) 
        (A => CO0) = (1.0, 1.0);
    if (B===1'b0 && NCI0===1'b0 && NCI1===1'b1) 
        (A => CO0) = (1.0, 1.0);
    if (B===1'b1 && NCI0===1'b1 && NCI1===1'b0) 
        (A => CO0) = (1.0, 1.0);
    if (B===1'b1 && NCI0===1'b1 && NCI1===1'b1) 
        (A => CO0) = (1.0, 1.0);
    ifnone
        (A => CO0) = (1.0, 1.0);

    // arc A --> CO1
    if (B===1'b0 && NCI0===1'b0 && NCI1===1'b0) 
        (A => CO1) = (1.0, 1.0);
    if (B===1'b0 && NCI0===1'b1 && NCI1===1'b0) 
        (A => CO1) = (1.0, 1.0);
    if (B===1'b1 && NCI0===1'b0 && NCI1===1'b1) 
        (A => CO1) = (1.0, 1.0);
    if (B===1'b1 && NCI0===1'b1 && NCI1===1'b1) 
        (A => CO1) = (1.0, 1.0);
    ifnone
        (A => CO1) = (1.0, 1.0);

    // arc B --> CO0
    if (A===1'b0 && NCI0===1'b0 && NCI1===1'b0) 
        (B => CO0) = (1.0, 1.0);
    if (A===1'b0 && NCI0===1'b0 && NCI1===1'b1) 
        (B => CO0) = (1.0, 1.0);
    if (A===1'b1 && NCI0===1'b1 && NCI1===1'b0) 
        (B => CO0) = (1.0, 1.0);
    if (A===1'b1 && NCI0===1'b1 && NCI1===1'b1) 
        (B => CO0) = (1.0, 1.0);
    ifnone
        (B => CO0) = (1.0, 1.0);

    // arc B --> CO1
    if (A===1'b0 && NCI0===1'b0 && NCI1===1'b0) 
        (B => CO1) = (1.0, 1.0);
    if (A===1'b0 && NCI0===1'b1 && NCI1===1'b0) 
        (B => CO1) = (1.0, 1.0);
    if (A===1'b1 && NCI0===1'b0 && NCI1===1'b1) 
        (B => CO1) = (1.0, 1.0);
    if (A===1'b1 && NCI0===1'b1 && NCI1===1'b1) 
        (B => CO1) = (1.0, 1.0);
    ifnone
        (B => CO1) = (1.0, 1.0);

    // arc NCI0 --> CO0
    if (A===1'b0 && B===1'b1 && NCI1===1'b0) 
        (NCI0 => CO0) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && NCI1===1'b1) 
        (NCI0 => CO0) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && NCI1===1'b0) 
        (NCI0 => CO0) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && NCI1===1'b1) 
        (NCI0 => CO0) = (1.0, 1.0);
    ifnone
        (NCI0 => CO0) = (1.0, 1.0);

    // arc NCI1 --> CO1
    if (A===1'b0 && B===1'b1 && NCI0===1'b0) 
        (NCI1 => CO1) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && NCI0===1'b1) 
        (NCI1 => CO1) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && NCI0===1'b0) 
        (NCI1 => CO1) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && NCI0===1'b1) 
        (NCI1 => CO1) = (1.0, 1.0);
    ifnone
        (NCI1 => CO1) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ADCSCM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:03:31 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module ADCSCM4N ( CO0, CO1, A, B, NCI0, NCI1 );
   input A, B, NCI0, NCI1;
   output CO0, CO1;
      ADCSCM2N_UDP4(CO0, A, B, NCI0);
      ADCSCM2N_UDP5(CO1, A, B, NCI1);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO0
    if (B===1'b0 && NCI0===1'b0 && NCI1===1'b0) 
        (A => CO0) = (1.0, 1.0);
    if (B===1'b0 && NCI0===1'b0 && NCI1===1'b1) 
        (A => CO0) = (1.0, 1.0);
    if (B===1'b1 && NCI0===1'b1 && NCI1===1'b0) 
        (A => CO0) = (1.0, 1.0);
    if (B===1'b1 && NCI0===1'b1 && NCI1===1'b1) 
        (A => CO0) = (1.0, 1.0);
    ifnone
        (A => CO0) = (1.0, 1.0);

    // arc A --> CO1
    if (B===1'b0 && NCI0===1'b0 && NCI1===1'b0) 
        (A => CO1) = (1.0, 1.0);
    if (B===1'b0 && NCI0===1'b1 && NCI1===1'b0) 
        (A => CO1) = (1.0, 1.0);
    if (B===1'b1 && NCI0===1'b0 && NCI1===1'b1) 
        (A => CO1) = (1.0, 1.0);
    if (B===1'b1 && NCI0===1'b1 && NCI1===1'b1) 
        (A => CO1) = (1.0, 1.0);
    ifnone
        (A => CO1) = (1.0, 1.0);

    // arc B --> CO0
    if (A===1'b0 && NCI0===1'b0 && NCI1===1'b0) 
        (B => CO0) = (1.0, 1.0);
    if (A===1'b0 && NCI0===1'b0 && NCI1===1'b1) 
        (B => CO0) = (1.0, 1.0);
    if (A===1'b1 && NCI0===1'b1 && NCI1===1'b0) 
        (B => CO0) = (1.0, 1.0);
    if (A===1'b1 && NCI0===1'b1 && NCI1===1'b1) 
        (B => CO0) = (1.0, 1.0);
    ifnone
        (B => CO0) = (1.0, 1.0);

    // arc B --> CO1
    if (A===1'b0 && NCI0===1'b0 && NCI1===1'b0) 
        (B => CO1) = (1.0, 1.0);
    if (A===1'b0 && NCI0===1'b1 && NCI1===1'b0) 
        (B => CO1) = (1.0, 1.0);
    if (A===1'b1 && NCI0===1'b0 && NCI1===1'b1) 
        (B => CO1) = (1.0, 1.0);
    if (A===1'b1 && NCI0===1'b1 && NCI1===1'b1) 
        (B => CO1) = (1.0, 1.0);
    ifnone
        (B => CO1) = (1.0, 1.0);

    // arc NCI0 --> CO0
    if (A===1'b0 && B===1'b1 && NCI1===1'b0) 
        (NCI0 => CO0) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && NCI1===1'b1) 
        (NCI0 => CO0) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && NCI1===1'b0) 
        (NCI0 => CO0) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && NCI1===1'b1) 
        (NCI0 => CO0) = (1.0, 1.0);
    ifnone
        (NCI0 => CO0) = (1.0, 1.0);

    // arc NCI1 --> CO1
    if (A===1'b0 && B===1'b1 && NCI0===1'b0) 
        (NCI1 => CO1) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && NCI0===1'b1) 
        (NCI1 => CO1) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && NCI0===1'b0) 
        (NCI1 => CO1) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && NCI0===1'b1) 
        (NCI1 => CO1) = (1.0, 1.0);
    ifnone
        (NCI1 => CO1) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ADCSCM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:06:32 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADCSIOM2N(A, B, CO0B, CO1B);
  input A, B;
  output CO0B, CO1B;

    nand SMC_I0(CO0B, A, B);

    not SMC_I1(A_bar, A);
    not SMC_I2(B_bar, B);
    and SMC_I3(CO1B, A_bar, B_bar);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO0B
    (A => CO0B) = (1.0, 1.0);

    // arc A --> CO1B
    (A => CO1B) = (1.0, 1.0);

    // arc B --> CO0B
    (B => CO0B) = (1.0, 1.0);

    // arc B --> CO1B
    (B => CO1B) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ADCSIOM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:07:36 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADCSIOM4N(A, B, CO0B, CO1B);
  input A, B;
  output CO0B, CO1B;

    nand SMC_I0(CO0B, A, B);

    not SMC_I1(A_bar, A);
    not SMC_I2(B_bar, B);
    and SMC_I3(CO1B, A_bar, B_bar);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO0B
    (A => CO0B) = (1.0, 1.0);

    // arc A --> CO1B
    (A => CO1B) = (1.0, 1.0);

    // arc B --> CO0B
    (B => CO0B) = (1.0, 1.0);

    // arc B --> CO1B
    (B => CO1B) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ADCSIOM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:06:03 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module ADCSOM2N ( CO0B, CO1B, A, B, CI0, CI1 );
   input A, B, CI0, CI1;
   output CO0B, CO1B;
      ADCSOM2N_UDP4(CO0B, A, B, CI0);
      ADCSOM2N_UDP5(CO1B, A, B, CI1);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO0B
    if (B===1'b0 && CI0===1'b1 && CI1===1'b0) 
        (A => CO0B) = (1.0, 1.0);
    if (B===1'b0 && CI0===1'b1 && CI1===1'b1) 
        (A => CO0B) = (1.0, 1.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b0) 
        (A => CO0B) = (1.0, 1.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b1) 
        (A => CO0B) = (1.0, 1.0);
    ifnone
        (A => CO0B) = (1.0, 1.0);

    // arc A --> CO1B
    if (B===1'b0 && CI0===1'b0 && CI1===1'b1) 
        (A => CO1B) = (1.0, 1.0);
    if (B===1'b0 && CI0===1'b1 && CI1===1'b1) 
        (A => CO1B) = (1.0, 1.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b0) 
        (A => CO1B) = (1.0, 1.0);
    if (B===1'b1 && CI0===1'b1 && CI1===1'b0) 
        (A => CO1B) = (1.0, 1.0);
    ifnone
        (A => CO1B) = (1.0, 1.0);

    // arc B --> CO0B
    if (A===1'b0 && CI0===1'b1 && CI1===1'b0) 
        (B => CO0B) = (1.0, 1.0);
    if (A===1'b0 && CI0===1'b1 && CI1===1'b1) 
        (B => CO0B) = (1.0, 1.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b0) 
        (B => CO0B) = (1.0, 1.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b1) 
        (B => CO0B) = (1.0, 1.0);
    ifnone
        (B => CO0B) = (1.0, 1.0);

    // arc B --> CO1B
    if (A===1'b0 && CI0===1'b0 && CI1===1'b1) 
        (B => CO1B) = (1.0, 1.0);
    if (A===1'b0 && CI0===1'b1 && CI1===1'b1) 
        (B => CO1B) = (1.0, 1.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b0) 
        (B => CO1B) = (1.0, 1.0);
    if (A===1'b1 && CI0===1'b1 && CI1===1'b0) 
        (B => CO1B) = (1.0, 1.0);
    ifnone
        (B => CO1B) = (1.0, 1.0);

    // arc CI0 --> CO0B
    if (A===1'b0 && B===1'b1 && CI1===1'b0) 
        (CI0 => CO0B) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && CI1===1'b1) 
        (CI0 => CO0B) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CI1===1'b0) 
        (CI0 => CO0B) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CI1===1'b1) 
        (CI0 => CO0B) = (1.0, 1.0);
    ifnone
        (CI0 => CO0B) = (1.0, 1.0);

    // arc CI1 --> CO1B
    if (A===1'b0 && B===1'b1 && CI0===1'b0) 
        (CI1 => CO1B) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && CI0===1'b1) 
        (CI1 => CO1B) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CI0===1'b0) 
        (CI1 => CO1B) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CI0===1'b1) 
        (CI1 => CO1B) = (1.0, 1.0);
    ifnone
        (CI1 => CO1B) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ADCSOM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:01:19 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module ADCSOM4N ( CO0B, CO1B, A, B, CI0, CI1 );
   input A, B, CI0, CI1;
   output CO0B, CO1B;
      ADCSOM2N_UDP4(CO0B, A, B, CI0);
      ADCSOM2N_UDP5(CO1B, A, B, CI1);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO0B
    if (B===1'b0 && CI0===1'b1 && CI1===1'b0) 
        (A => CO0B) = (1.0, 1.0);
    if (B===1'b0 && CI0===1'b1 && CI1===1'b1) 
        (A => CO0B) = (1.0, 1.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b0) 
        (A => CO0B) = (1.0, 1.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b1) 
        (A => CO0B) = (1.0, 1.0);
    ifnone
        (A => CO0B) = (1.0, 1.0);

    // arc A --> CO1B
    if (B===1'b0 && CI0===1'b0 && CI1===1'b1) 
        (A => CO1B) = (1.0, 1.0);
    if (B===1'b0 && CI0===1'b1 && CI1===1'b1) 
        (A => CO1B) = (1.0, 1.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b0) 
        (A => CO1B) = (1.0, 1.0);
    if (B===1'b1 && CI0===1'b1 && CI1===1'b0) 
        (A => CO1B) = (1.0, 1.0);
    ifnone
        (A => CO1B) = (1.0, 1.0);

    // arc B --> CO0B
    if (A===1'b0 && CI0===1'b1 && CI1===1'b0) 
        (B => CO0B) = (1.0, 1.0);
    if (A===1'b0 && CI0===1'b1 && CI1===1'b1) 
        (B => CO0B) = (1.0, 1.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b0) 
        (B => CO0B) = (1.0, 1.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b1) 
        (B => CO0B) = (1.0, 1.0);
    ifnone
        (B => CO0B) = (1.0, 1.0);

    // arc B --> CO1B
    if (A===1'b0 && CI0===1'b0 && CI1===1'b1) 
        (B => CO1B) = (1.0, 1.0);
    if (A===1'b0 && CI0===1'b1 && CI1===1'b1) 
        (B => CO1B) = (1.0, 1.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b0) 
        (B => CO1B) = (1.0, 1.0);
    if (A===1'b1 && CI0===1'b1 && CI1===1'b0) 
        (B => CO1B) = (1.0, 1.0);
    ifnone
        (B => CO1B) = (1.0, 1.0);

    // arc CI0 --> CO0B
    if (A===1'b0 && B===1'b1 && CI1===1'b0) 
        (CI0 => CO0B) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && CI1===1'b1) 
        (CI0 => CO0B) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CI1===1'b0) 
        (CI0 => CO0B) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CI1===1'b1) 
        (CI0 => CO0B) = (1.0, 1.0);
    ifnone
        (CI0 => CO0B) = (1.0, 1.0);

    // arc CI1 --> CO1B
    if (A===1'b0 && B===1'b1 && CI0===1'b0) 
        (CI1 => CO1B) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && CI0===1'b1) 
        (CI1 => CO1B) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CI0===1'b0) 
        (CI1 => CO1B) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CI0===1'b1) 
        (CI1 => CO1B) = (1.0, 1.0);
    ifnone
        (CI1 => CO1B) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ADCSOM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:03:49 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module ADFCGCM2N ( CO, A, B, NCI );
   input A, B, NCI;
   output CO;
      ADFCGCM2N_UDP3(CO, A, B, NCI);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO
    if (B===1'b0 && NCI===1'b0) 
        (A => CO) = (1.0, 1.0);
    if (B===1'b1 && NCI===1'b1) 
        (A => CO) = (1.0, 1.0);
    ifnone
        (A => CO) = (1.0, 1.0);

    // arc B --> CO
    if (A===1'b0 && NCI===1'b0) 
        (B => CO) = (1.0, 1.0);
    if (A===1'b1 && NCI===1'b1) 
        (B => CO) = (1.0, 1.0);
    ifnone
        (B => CO) = (1.0, 1.0);

    // arc NCI --> CO
    if (A===1'b0 && B===1'b1) 
        (NCI => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0) 
        (NCI => CO) = (1.0, 1.0);
    ifnone
        (NCI => CO) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ADFCGCM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:06:34 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module ADFCGCM4N ( CO, A, B, NCI );
   input A, B, NCI;
   output CO;
      ADFCGCM2N_UDP3(CO, A, B, NCI);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO
    if (B===1'b0 && NCI===1'b0) 
        (A => CO) = (1.0, 1.0);
    if (B===1'b1 && NCI===1'b1) 
        (A => CO) = (1.0, 1.0);
    ifnone
        (A => CO) = (1.0, 1.0);

    // arc B --> CO
    if (A===1'b0 && NCI===1'b0) 
        (B => CO) = (1.0, 1.0);
    if (A===1'b1 && NCI===1'b1) 
        (B => CO) = (1.0, 1.0);
    ifnone
        (B => CO) = (1.0, 1.0);

    // arc NCI --> CO
    if (A===1'b0 && B===1'b1) 
        (NCI => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0) 
        (NCI => CO) = (1.0, 1.0);
    ifnone
        (NCI => CO) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ADFCGCM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:01:23 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module ADFCGOM2N ( COB, A, B, CI );
   input A, B, CI;
   output COB;
      ADFCGOM2N_UDP3(COB, A, B, CI);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> COB
    if (B===1'b0 && CI===1'b1) 
        (A => COB) = (1.0, 1.0);
    if (B===1'b1 && CI===1'b0) 
        (A => COB) = (1.0, 1.0);
    ifnone
        (A => COB) = (1.0, 1.0);

    // arc B --> COB
    if (A===1'b0 && CI===1'b1) 
        (B => COB) = (1.0, 1.0);
    if (A===1'b1 && CI===1'b0) 
        (B => COB) = (1.0, 1.0);
    ifnone
        (B => COB) = (1.0, 1.0);

    // arc CI --> COB
    if (A===1'b0 && B===1'b1) 
        (CI => COB) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0) 
        (CI => COB) = (1.0, 1.0);
    ifnone
        (CI => COB) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ADFCGOM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:06:07 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module ADFCGOM4N ( COB, A, B, CI );
   input A, B, CI;
   output COB;
      ADFCGOM2N_UDP3(COB, A, B, CI);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> COB
    if (B===1'b0 && CI===1'b1) 
        (A => COB) = (1.0, 1.0);
    if (B===1'b1 && CI===1'b0) 
        (A => COB) = (1.0, 1.0);
    ifnone
        (A => COB) = (1.0, 1.0);

    // arc B --> COB
    if (A===1'b0 && CI===1'b1) 
        (B => COB) = (1.0, 1.0);
    if (A===1'b1 && CI===1'b0) 
        (B => COB) = (1.0, 1.0);
    ifnone
        (B => COB) = (1.0, 1.0);

    // arc CI --> COB
    if (A===1'b0 && B===1'b1) 
        (CI => COB) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0) 
        (CI => COB) = (1.0, 1.0);
    ifnone
        (CI => COB) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ADFCGOM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:03:55 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module ADFCM2N ( CO, S, A, B, NCI );
   input A, B, NCI;
   output CO, S;
      ADFCM2N_UDP3(CO, A, B, NCI);
      ADFCM2N_UDP4(S, A, B, NCI);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO
    if (B===1'b0 && NCI===1'b0) 
        (A => CO) = (1.0, 1.0);
    if (B===1'b1 && NCI===1'b1) 
        (A => CO) = (1.0, 1.0);
    ifnone
        (A => CO) = (1.0, 1.0);

    // arc A --> S
    if (B===1'b0 && NCI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && NCI===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && NCI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && NCI===1'b1) 
        (A => S) = (1.0, 1.0);
    ifnone
        ( posedge A => ( S +: A ) ) = (1.0, 1.0);
        ( negedge A => ( S +: A ) ) = (1.0, 1.0);

    // arc B --> CO
    if (A===1'b0 && NCI===1'b0) 
        (B => CO) = (1.0, 1.0);
    if (A===1'b1 && NCI===1'b1) 
        (B => CO) = (1.0, 1.0);
    ifnone
        (B => CO) = (1.0, 1.0);

    // arc B --> S
    if (A===1'b0 && NCI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && NCI===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && NCI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && NCI===1'b1) 
        (B => S) = (1.0, 1.0);
    ifnone
        ( posedge B => ( S +: B ) ) = (1.0, 1.0);
        ( negedge B => ( S +: B ) ) = (1.0, 1.0);

    // arc NCI --> CO
    if (A===1'b0 && B===1'b1) 
        (NCI => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0) 
        (NCI => CO) = (1.0, 1.0);
    ifnone
        (NCI => CO) = (1.0, 1.0);

    // arc NCI --> S
    if (A===1'b0 && B===1'b0) 
        (NCI => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1) 
        (NCI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0) 
        (NCI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1) 
        (NCI => S) = (1.0, 1.0);
    ifnone
        ( posedge NCI => ( S +: NCI ) ) = (1.0, 1.0);
        ( negedge NCI => ( S +: NCI ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ADFCM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:03:32 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module ADFCM4N ( CO, S, A, B, NCI );
   input A, B, NCI;
   output CO, S;
      ADFCM2N_UDP3(CO, A, B, NCI);
      ADFCM2N_UDP4(S, A, B, NCI);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO
    if (B===1'b0 && NCI===1'b0) 
        (A => CO) = (1.0, 1.0);
    if (B===1'b1 && NCI===1'b1) 
        (A => CO) = (1.0, 1.0);
    ifnone
        (A => CO) = (1.0, 1.0);

    // arc A --> S
    if (B===1'b0 && NCI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && NCI===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && NCI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && NCI===1'b1) 
        (A => S) = (1.0, 1.0);
    ifnone
        ( posedge A => ( S +: A ) ) = (1.0, 1.0);
        ( negedge A => ( S +: A ) ) = (1.0, 1.0);

    // arc B --> CO
    if (A===1'b0 && NCI===1'b0) 
        (B => CO) = (1.0, 1.0);
    if (A===1'b1 && NCI===1'b1) 
        (B => CO) = (1.0, 1.0);
    ifnone
        (B => CO) = (1.0, 1.0);

    // arc B --> S
    if (A===1'b0 && NCI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && NCI===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && NCI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && NCI===1'b1) 
        (B => S) = (1.0, 1.0);
    ifnone
        ( posedge B => ( S +: B ) ) = (1.0, 1.0);
        ( negedge B => ( S +: B ) ) = (1.0, 1.0);

    // arc NCI --> CO
    if (A===1'b0 && B===1'b1) 
        (NCI => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0) 
        (NCI => CO) = (1.0, 1.0);
    ifnone
        (NCI => CO) = (1.0, 1.0);

    // arc NCI --> S
    if (A===1'b0 && B===1'b0) 
        (NCI => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1) 
        (NCI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0) 
        (NCI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1) 
        (NCI => S) = (1.0, 1.0);
    ifnone
        ( posedge NCI => ( S +: NCI ) ) = (1.0, 1.0);
        ( negedge NCI => ( S +: NCI ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ADFCM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:08:36 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module ADFCSCM2N ( CO0, CO1, S, A, B, CS, NCI0, NCI1 );
   input A, B, CS, NCI0, NCI1;
   output CO0, CO1, S;
      ADFCSCM2N_UDP5(CO0, A, B, NCI0);
      ADFCSCM2N_UDP6(CO1, A, B, NCI1);
      ADFCSCM2N_UDP7(S, A, B, CS, NCI0, NCI1);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO0
    if (B===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0) 
        (A => CO0) = (1.0, 1.0);
    if (B===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1) 
        (A => CO0) = (1.0, 1.0);
    if (B===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0) 
        (A => CO0) = (1.0, 1.0);
    if (B===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1) 
        (A => CO0) = (1.0, 1.0);
    if (B===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0) 
        (A => CO0) = (1.0, 1.0);
    if (B===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1) 
        (A => CO0) = (1.0, 1.0);
    if (B===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0) 
        (A => CO0) = (1.0, 1.0);
    if (B===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1) 
        (A => CO0) = (1.0, 1.0);
    ifnone
        (A => CO0) = (1.0, 1.0);

    // arc A --> CO1
    if (B===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0) 
        (A => CO1) = (1.0, 1.0);
    if (B===1'b0 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0) 
        (A => CO1) = (1.0, 1.0);
    if (B===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0) 
        (A => CO1) = (1.0, 1.0);
    if (B===1'b0 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0) 
        (A => CO1) = (1.0, 1.0);
    if (B===1'b1 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1) 
        (A => CO1) = (1.0, 1.0);
    if (B===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1) 
        (A => CO1) = (1.0, 1.0);
    if (B===1'b1 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1) 
        (A => CO1) = (1.0, 1.0);
    if (B===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1) 
        (A => CO1) = (1.0, 1.0);
    ifnone
        (A => CO1) = (1.0, 1.0);

    // arc A --> S
    if (B===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1) 
        (A => S) = (1.0, 1.0);
    ifnone
        ( posedge A => ( S +: A ) ) = (1.0, 1.0);
        ( negedge A => ( S +: A ) ) = (1.0, 1.0);

    // arc B --> CO0
    if (A===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0) 
        (B => CO0) = (1.0, 1.0);
    if (A===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1) 
        (B => CO0) = (1.0, 1.0);
    if (A===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0) 
        (B => CO0) = (1.0, 1.0);
    if (A===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1) 
        (B => CO0) = (1.0, 1.0);
    if (A===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0) 
        (B => CO0) = (1.0, 1.0);
    if (A===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1) 
        (B => CO0) = (1.0, 1.0);
    if (A===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0) 
        (B => CO0) = (1.0, 1.0);
    if (A===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1) 
        (B => CO0) = (1.0, 1.0);
    ifnone
        (B => CO0) = (1.0, 1.0);

    // arc B --> CO1
    if (A===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0) 
        (B => CO1) = (1.0, 1.0);
    if (A===1'b0 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0) 
        (B => CO1) = (1.0, 1.0);
    if (A===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0) 
        (B => CO1) = (1.0, 1.0);
    if (A===1'b0 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0) 
        (B => CO1) = (1.0, 1.0);
    if (A===1'b1 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1) 
        (B => CO1) = (1.0, 1.0);
    if (A===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1) 
        (B => CO1) = (1.0, 1.0);
    if (A===1'b1 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1) 
        (B => CO1) = (1.0, 1.0);
    if (A===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1) 
        (B => CO1) = (1.0, 1.0);
    ifnone
        (B => CO1) = (1.0, 1.0);

    // arc B --> S
    if (A===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1) 
        (B => S) = (1.0, 1.0);
    ifnone
        ( posedge B => ( S +: B ) ) = (1.0, 1.0);
        ( negedge B => ( S +: B ) ) = (1.0, 1.0);

    // arc CS --> S
    if (A===1'b0 && B===1'b0 && NCI0===1'b0 && NCI1===1'b1) 
        (CS => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && NCI0===1'b1 && NCI1===1'b0) 
        (CS => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && NCI0===1'b0 && NCI1===1'b1) 
        (CS => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && NCI0===1'b1 && NCI1===1'b0) 
        (CS => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && NCI0===1'b0 && NCI1===1'b1) 
        (CS => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && NCI0===1'b1 && NCI1===1'b0) 
        (CS => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && NCI0===1'b0 && NCI1===1'b1) 
        (CS => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && NCI0===1'b1 && NCI1===1'b0) 
        (CS => S) = (1.0, 1.0);
    ifnone
        ( posedge CS => ( S +: CS ) ) = (1.0, 1.0);
        ( negedge CS => ( S +: CS ) ) = (1.0, 1.0);

    // arc NCI0 --> CO0
    if (A===1'b0 && B===1'b1 && CS===1'b0 && NCI1===1'b0) 
        (NCI0 => CO0) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && CS===1'b0 && NCI1===1'b1) 
        (NCI0 => CO0) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && CS===1'b1 && NCI1===1'b0) 
        (NCI0 => CO0) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && CS===1'b1 && NCI1===1'b1) 
        (NCI0 => CO0) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CS===1'b0 && NCI1===1'b0) 
        (NCI0 => CO0) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CS===1'b0 && NCI1===1'b1) 
        (NCI0 => CO0) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CS===1'b1 && NCI1===1'b0) 
        (NCI0 => CO0) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CS===1'b1 && NCI1===1'b1) 
        (NCI0 => CO0) = (1.0, 1.0);
    ifnone
        (NCI0 => CO0) = (1.0, 1.0);

    // arc NCI0 --> S
    if (A===1'b0 && B===1'b0 && NCI1===1'b0) 
        (NCI0 => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && NCI1===1'b1) 
        (NCI0 => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && NCI1===1'b0) 
        (NCI0 => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && NCI1===1'b1) 
        (NCI0 => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && NCI1===1'b0) 
        (NCI0 => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && NCI1===1'b1) 
        (NCI0 => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && NCI1===1'b0) 
        (NCI0 => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && NCI1===1'b1) 
        (NCI0 => S) = (1.0, 1.0);
    ifnone
        ( posedge NCI0 => ( S +: NCI0 ) ) = (1.0, 1.0);
        ( negedge NCI0 => ( S +: NCI0 ) ) = (1.0, 1.0);

    // arc NCI1 --> CO1
    if (A===1'b0 && B===1'b1 && CS===1'b0 && NCI0===1'b0) 
        (NCI1 => CO1) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && CS===1'b0 && NCI0===1'b1) 
        (NCI1 => CO1) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && CS===1'b1 && NCI0===1'b0) 
        (NCI1 => CO1) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && CS===1'b1 && NCI0===1'b1) 
        (NCI1 => CO1) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CS===1'b0 && NCI0===1'b0) 
        (NCI1 => CO1) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CS===1'b0 && NCI0===1'b1) 
        (NCI1 => CO1) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CS===1'b1 && NCI0===1'b0) 
        (NCI1 => CO1) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CS===1'b1 && NCI0===1'b1) 
        (NCI1 => CO1) = (1.0, 1.0);
    ifnone
        (NCI1 => CO1) = (1.0, 1.0);

    // arc NCI1 --> S
    if (A===1'b0 && B===1'b0 && NCI0===1'b0) 
        (NCI1 => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && NCI0===1'b1) 
        (NCI1 => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && NCI0===1'b0) 
        (NCI1 => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && NCI0===1'b1) 
        (NCI1 => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && NCI0===1'b0) 
        (NCI1 => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && NCI0===1'b1) 
        (NCI1 => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && NCI0===1'b0) 
        (NCI1 => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && NCI0===1'b1) 
        (NCI1 => S) = (1.0, 1.0);
    ifnone
        ( posedge NCI1 => ( S +: NCI1 ) ) = (1.0, 1.0);
        ( negedge NCI1 => ( S +: NCI1 ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ADFCSCM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:07:35 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module ADFCSCM4N ( CO0, CO1, S, A, B, CS, NCI0, NCI1 );
   input A, B, CS, NCI0, NCI1;
   output CO0, CO1, S;
      ADFCSCM2N_UDP5(CO0, A, B, NCI0);
      ADFCSCM2N_UDP6(CO1, A, B, NCI1);
      ADFCSCM2N_UDP7(S, A, B, CS, NCI0, NCI1);
   
  `ifdef functional // functional //

  `else // functional //

 specify


    // arc A --> CO0
    if (B===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0) 
        (A => CO0) = (1.0, 1.0);
    if (B===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1) 
        (A => CO0) = (1.0, 1.0);
    if (B===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0) 
        (A => CO0) = (1.0, 1.0);
    if (B===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1) 
        (A => CO0) = (1.0, 1.0);
    if (B===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0) 
        (A => CO0) = (1.0, 1.0);
    if (B===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1) 
        (A => CO0) = (1.0, 1.0);
    if (B===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0) 
        (A => CO0) = (1.0, 1.0);
    if (B===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1) 
        (A => CO0) = (1.0, 1.0);
    ifnone
        (A => CO0) = (1.0, 1.0);

    // arc A --> CO1
    if (B===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0) 
        (A => CO1) = (1.0, 1.0);
    if (B===1'b0 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0) 
        (A => CO1) = (1.0, 1.0);
    if (B===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0) 
        (A => CO1) = (1.0, 1.0);
    if (B===1'b0 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0) 
        (A => CO1) = (1.0, 1.0);
    if (B===1'b1 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1) 
        (A => CO1) = (1.0, 1.0);
    if (B===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1) 
        (A => CO1) = (1.0, 1.0);
    if (B===1'b1 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1) 
        (A => CO1) = (1.0, 1.0);
    if (B===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1) 
        (A => CO1) = (1.0, 1.0);
    ifnone
        (A => CO1) = (1.0, 1.0);

    // arc A --> S
    if (B===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1) 
        (A => S) = (1.0, 1.0);
    ifnone
        ( posedge A => ( S +: A ) ) = (1.0, 1.0);
        ( negedge A => ( S +: A ) ) = (1.0, 1.0);

    // arc B --> CO0
    if (A===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0) 
        (B => CO0) = (1.0, 1.0);
    if (A===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1) 
        (B => CO0) = (1.0, 1.0);
    if (A===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0) 
        (B => CO0) = (1.0, 1.0);
    if (A===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1) 
        (B => CO0) = (1.0, 1.0);
    if (A===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0) 
        (B => CO0) = (1.0, 1.0);
    if (A===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1) 
        (B => CO0) = (1.0, 1.0);
    if (A===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0) 
        (B => CO0) = (1.0, 1.0);
    if (A===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1) 
        (B => CO0) = (1.0, 1.0);
    ifnone
        (B => CO0) = (1.0, 1.0);

    // arc B --> CO1
    if (A===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0) 
        (B => CO1) = (1.0, 1.0);
    if (A===1'b0 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0) 
        (B => CO1) = (1.0, 1.0);
    if (A===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0) 
        (B => CO1) = (1.0, 1.0);
    if (A===1'b0 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0) 
        (B => CO1) = (1.0, 1.0);
    if (A===1'b1 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1) 
        (B => CO1) = (1.0, 1.0);
    if (A===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1) 
        (B => CO1) = (1.0, 1.0);
    if (A===1'b1 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1) 
        (B => CO1) = (1.0, 1.0);
    if (A===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1) 
        (B => CO1) = (1.0, 1.0);
    ifnone
        (B => CO1) = (1.0, 1.0);

    // arc B --> S
    if (A===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1) 
        (B => S) = (1.0, 1.0);
    ifnone
        ( posedge B => ( S +: B ) ) = (1.0, 1.0);
        ( negedge B => ( S +: B ) ) = (1.0, 1.0);

    // arc CS --> S
    if (A===1'b0 && B===1'b0 && NCI0===1'b0 && NCI1===1'b1) 
        (CS => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && NCI0===1'b1 && NCI1===1'b0) 
        (CS => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && NCI0===1'b0 && NCI1===1'b1) 
        (CS => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && NCI0===1'b1 && NCI1===1'b0) 
        (CS => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && NCI0===1'b0 && NCI1===1'b1) 
        (CS => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && NCI0===1'b1 && NCI1===1'b0) 
        (CS => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && NCI0===1'b0 && NCI1===1'b1) 
        (CS => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && NCI0===1'b1 && NCI1===1'b0) 
        (CS => S) = (1.0, 1.0);
    ifnone
        ( posedge CS => ( S +: CS ) ) = (1.0, 1.0);
        ( negedge CS => ( S +: CS ) ) = (1.0, 1.0);

    // arc NCI0 --> CO0
    if (A===1'b0 && B===1'b1 && CS===1'b0 && NCI1===1'b0) 
        (NCI0 => CO0) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && CS===1'b0 && NCI1===1'b1) 
        (NCI0 => CO0) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && CS===1'b1 && NCI1===1'b0) 
        (NCI0 => CO0) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && CS===1'b1 && NCI1===1'b1) 
        (NCI0 => CO0) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CS===1'b0 && NCI1===1'b0) 
        (NCI0 => CO0) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CS===1'b0 && NCI1===1'b1) 
        (NCI0 => CO0) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CS===1'b1 && NCI1===1'b0) 
        (NCI0 => CO0) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CS===1'b1 && NCI1===1'b1) 
        (NCI0 => CO0) = (1.0, 1.0);
    ifnone
        (NCI0 => CO0) = (1.0, 1.0);

    // arc NCI0 --> S
    if (A===1'b0 && B===1'b0 && NCI1===1'b0) 
        (NCI0 => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && NCI1===1'b1) 
        (NCI0 => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && NCI1===1'b0) 
        (NCI0 => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && NCI1===1'b1) 
        (NCI0 => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && NCI1===1'b0) 
        (NCI0 => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && NCI1===1'b1) 
        (NCI0 => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && NCI1===1'b0) 
        (NCI0 => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && NCI1===1'b1) 
        (NCI0 => S) = (1.0, 1.0);
    ifnone
        ( posedge NCI0 => ( S +: NCI0 ) ) = (1.0, 1.0);
        ( negedge NCI0 => ( S +: NCI0 ) ) = (1.0, 1.0);

    // arc NCI1 --> CO1
    if (A===1'b0 && B===1'b1 && CS===1'b0 && NCI0===1'b0) 
        (NCI1 => CO1) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && CS===1'b0 && NCI0===1'b1) 
        (NCI1 => CO1) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && CS===1'b1 && NCI0===1'b0) 
        (NCI1 => CO1) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && CS===1'b1 && NCI0===1'b1) 
        (NCI1 => CO1) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CS===1'b0 && NCI0===1'b0) 
        (NCI1 => CO1) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CS===1'b0 && NCI0===1'b1) 
        (NCI1 => CO1) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CS===1'b1 && NCI0===1'b0) 
        (NCI1 => CO1) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CS===1'b1 && NCI0===1'b1) 
        (NCI1 => CO1) = (1.0, 1.0);
    ifnone
        (NCI1 => CO1) = (1.0, 1.0);

    // arc NCI1 --> S
    if (A===1'b0 && B===1'b0 && NCI0===1'b0) 
        (NCI1 => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && NCI0===1'b1) 
        (NCI1 => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && NCI0===1'b0) 
        (NCI1 => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && NCI0===1'b1) 
        (NCI1 => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && NCI0===1'b0) 
        (NCI1 => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && NCI0===1'b1) 
        (NCI1 => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && NCI0===1'b0) 
        (NCI1 => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && NCI0===1'b1) 
        (NCI1 => S) = (1.0, 1.0);
    ifnone
        ( posedge NCI1 => ( S +: NCI1 ) ) = (1.0, 1.0);
        ( negedge NCI1 => ( S +: NCI1 ) ) = (1.0, 1.0);




  endspecify

  `endif // functional //
endmodule     // ADFCSCM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:06:05 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADFCSIOM2N(A, B, CS, CO0B, CO1B, S);
  input A, B, CS;
  output CO0B, CO1B, S;

    nand SMC_I0(CO0B, A, B);

    not SMC_I1(A_bar, A);
    not SMC_I2(B_bar, B);
    and SMC_I3(CO1B, A_bar, B_bar);

    xor SMC_I4(S, A, B, CS);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO0B
    if (CS===1'b0) 
        (A => CO0B) = (1.0, 1.0);
    if (CS===1'b1) 
        (A => CO0B) = (1.0, 1.0);
    ifnone
        (A => CO0B) = (1.0, 1.0);

    // arc A --> CO1B
    if (CS===1'b0) 
        (A => CO1B) = (1.0, 1.0);
    if (CS===1'b1) 
        (A => CO1B) = (1.0, 1.0);
    ifnone
        (A => CO1B) = (1.0, 1.0);

    // arc A --> S
    if (B===1'b0 && CS===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && CS===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CS===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CS===1'b1) 
        (A => S) = (1.0, 1.0);
    ifnone
        ( posedge A => ( S +: A ) ) = (1.0, 1.0);
        ( negedge A => ( S +: A ) ) = (1.0, 1.0);

    // arc B --> CO0B
    if (CS===1'b0) 
        (B => CO0B) = (1.0, 1.0);
    if (CS===1'b1) 
        (B => CO0B) = (1.0, 1.0);
    ifnone
        (B => CO0B) = (1.0, 1.0);

    // arc B --> CO1B
    if (CS===1'b0) 
        (B => CO1B) = (1.0, 1.0);
    if (CS===1'b1) 
        (B => CO1B) = (1.0, 1.0);
    ifnone
        (B => CO1B) = (1.0, 1.0);

    // arc B --> S
    if (A===1'b0 && CS===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && CS===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CS===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CS===1'b1) 
        (B => S) = (1.0, 1.0);
    ifnone
        ( posedge B => ( S +: B ) ) = (1.0, 1.0);
        ( negedge B => ( S +: B ) ) = (1.0, 1.0);

    // arc CS --> S
    if (A===1'b0 && B===1'b0) 
        (CS => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1) 
        (CS => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0) 
        (CS => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1) 
        (CS => S) = (1.0, 1.0);
    ifnone
        ( posedge CS => ( S +: CS ) ) = (1.0, 1.0);
        ( negedge CS => ( S +: CS ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ADFCSIOM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:02:49 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADFCSIOM4N(A, B, CS, CO0B, CO1B, S);
  input A, B, CS;
  output CO0B, CO1B, S;

    nand SMC_I0(CO0B, A, B);

    not SMC_I1(A_bar, A);
    not SMC_I2(B_bar, B);
    and SMC_I3(CO1B, A_bar, B_bar);

    xor SMC_I4(S, A, B, CS);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO0B
    if (CS===1'b0) 
        (A => CO0B) = (1.0, 1.0);
    if (CS===1'b1) 
        (A => CO0B) = (1.0, 1.0);
    ifnone
        (A => CO0B) = (1.0, 1.0);

    // arc A --> CO1B
    if (CS===1'b0) 
        (A => CO1B) = (1.0, 1.0);
    if (CS===1'b1) 
        (A => CO1B) = (1.0, 1.0);
    ifnone
        (A => CO1B) = (1.0, 1.0);

    // arc A --> S
    if (B===1'b0 && CS===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && CS===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CS===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CS===1'b1) 
        (A => S) = (1.0, 1.0);
    ifnone
        ( posedge A => ( S +: A ) ) = (1.0, 1.0);
        ( negedge A => ( S +: A ) ) = (1.0, 1.0);

    // arc B --> CO0B
    if (CS===1'b0) 
        (B => CO0B) = (1.0, 1.0);
    if (CS===1'b1) 
        (B => CO0B) = (1.0, 1.0);
    ifnone
        (B => CO0B) = (1.0, 1.0);

    // arc B --> CO1B
    if (CS===1'b0) 
        (B => CO1B) = (1.0, 1.0);
    if (CS===1'b1) 
        (B => CO1B) = (1.0, 1.0);
    ifnone
        (B => CO1B) = (1.0, 1.0);

    // arc B --> S
    if (A===1'b0 && CS===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && CS===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CS===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CS===1'b1) 
        (B => S) = (1.0, 1.0);
    ifnone
        ( posedge B => ( S +: B ) ) = (1.0, 1.0);
        ( negedge B => ( S +: B ) ) = (1.0, 1.0);

    // arc CS --> S
    if (A===1'b0 && B===1'b0) 
        (CS => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1) 
        (CS => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0) 
        (CS => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1) 
        (CS => S) = (1.0, 1.0);
    ifnone
        ( posedge CS => ( S +: CS ) ) = (1.0, 1.0);
        ( negedge CS => ( S +: CS ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ADFCSIOM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:07:15 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module ADFCSOM2N ( CO0B, CO1B, S, A, B, CI0, CI1, CS );
   input A, B, CI0, CI1, CS;
   output CO0B, CO1B, S;
      ADFCSOM2N_UDP5(CO0B, A, B, CI0);
      ADFCSOM2N_UDP6(CO1B, A, B, CI1);
      ADFCSOM2N_UDP7(S, A, B, CI0, CI1, CS);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO0B
    if (B===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b0) 
        (A => CO0B) = (1.0, 1.0);
    if (B===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b1) 
        (A => CO0B) = (1.0, 1.0);
    if (B===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b0) 
        (A => CO0B) = (1.0, 1.0);
    if (B===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b1) 
        (A => CO0B) = (1.0, 1.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b0) 
        (A => CO0B) = (1.0, 1.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b1) 
        (A => CO0B) = (1.0, 1.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b0) 
        (A => CO0B) = (1.0, 1.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b1) 
        (A => CO0B) = (1.0, 1.0);
    ifnone
        (A => CO0B) = (1.0, 1.0);

    // arc A --> CO1B
    if (B===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b0) 
        (A => CO1B) = (1.0, 1.0);
    if (B===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b1) 
        (A => CO1B) = (1.0, 1.0);
    if (B===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b0) 
        (A => CO1B) = (1.0, 1.0);
    if (B===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b1) 
        (A => CO1B) = (1.0, 1.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b0) 
        (A => CO1B) = (1.0, 1.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b1) 
        (A => CO1B) = (1.0, 1.0);
    if (B===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b0) 
        (A => CO1B) = (1.0, 1.0);
    if (B===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b1) 
        (A => CO1B) = (1.0, 1.0);
    ifnone
        (A => CO1B) = (1.0, 1.0);

    // arc A --> S
    if (B===1'b0 && CI0===1'b0 && CI1===1'b0 && CS===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && CI0===1'b0 && CI1===1'b0 && CS===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CI0===1'b1 && CI1===1'b1 && CS===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CI0===1'b1 && CI1===1'b1 && CS===1'b1) 
        (A => S) = (1.0, 1.0);
    ifnone
        ( posedge A => ( S +: A ) ) = (1.0, 1.0);
        ( negedge A => ( S +: A ) ) = (1.0, 1.0);

    // arc B --> CO0B
    if (A===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b0) 
        (B => CO0B) = (1.0, 1.0);
    if (A===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b1) 
        (B => CO0B) = (1.0, 1.0);
    if (A===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b0) 
        (B => CO0B) = (1.0, 1.0);
    if (A===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b1) 
        (B => CO0B) = (1.0, 1.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b0) 
        (B => CO0B) = (1.0, 1.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b1) 
        (B => CO0B) = (1.0, 1.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b0) 
        (B => CO0B) = (1.0, 1.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b1) 
        (B => CO0B) = (1.0, 1.0);
    ifnone
        (B => CO0B) = (1.0, 1.0);

    // arc B --> CO1B
    if (A===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b0) 
        (B => CO1B) = (1.0, 1.0);
    if (A===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b1) 
        (B => CO1B) = (1.0, 1.0);
    if (A===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b0) 
        (B => CO1B) = (1.0, 1.0);
    if (A===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b1) 
        (B => CO1B) = (1.0, 1.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b0) 
        (B => CO1B) = (1.0, 1.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b1) 
        (B => CO1B) = (1.0, 1.0);
    if (A===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b0) 
        (B => CO1B) = (1.0, 1.0);
    if (A===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b1) 
        (B => CO1B) = (1.0, 1.0);
    ifnone
        (B => CO1B) = (1.0, 1.0);

    // arc B --> S
    if (A===1'b0 && CI0===1'b0 && CI1===1'b0 && CS===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && CI0===1'b0 && CI1===1'b0 && CS===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CI0===1'b1 && CI1===1'b1 && CS===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CI0===1'b1 && CI1===1'b1 && CS===1'b1) 
        (B => S) = (1.0, 1.0);
    ifnone
        ( posedge B => ( S +: B ) ) = (1.0, 1.0);
        ( negedge B => ( S +: B ) ) = (1.0, 1.0);

    // arc CI0 --> CO0B
    if (A===1'b0 && B===1'b1 && CI1===1'b0 && CS===1'b0) 
        (CI0 => CO0B) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && CI1===1'b0 && CS===1'b1) 
        (CI0 => CO0B) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && CI1===1'b1 && CS===1'b0) 
        (CI0 => CO0B) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && CI1===1'b1 && CS===1'b1) 
        (CI0 => CO0B) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CI1===1'b0 && CS===1'b0) 
        (CI0 => CO0B) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CI1===1'b0 && CS===1'b1) 
        (CI0 => CO0B) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CI1===1'b1 && CS===1'b0) 
        (CI0 => CO0B) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CI1===1'b1 && CS===1'b1) 
        (CI0 => CO0B) = (1.0, 1.0);
    ifnone
        (CI0 => CO0B) = (1.0, 1.0);

    // arc CI0 --> S
    if (A===1'b0 && B===1'b0 && CI1===1'b0) 
        (CI0 => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && CI1===1'b1) 
        (CI0 => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && CI1===1'b0) 
        (CI0 => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && CI1===1'b1) 
        (CI0 => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CI1===1'b0) 
        (CI0 => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CI1===1'b1) 
        (CI0 => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && CI1===1'b0) 
        (CI0 => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && CI1===1'b1) 
        (CI0 => S) = (1.0, 1.0);
    ifnone
        ( posedge CI0 => ( S +: CI0 ) ) = (1.0, 1.0);
        ( negedge CI0 => ( S +: CI0 ) ) = (1.0, 1.0);

    // arc CI1 --> CO1B
    if (A===1'b0 && B===1'b1 && CI0===1'b0 && CS===1'b0) 
        (CI1 => CO1B) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && CI0===1'b0 && CS===1'b1) 
        (CI1 => CO1B) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && CI0===1'b1 && CS===1'b0) 
        (CI1 => CO1B) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && CI0===1'b1 && CS===1'b1) 
        (CI1 => CO1B) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CI0===1'b0 && CS===1'b0) 
        (CI1 => CO1B) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CI0===1'b0 && CS===1'b1) 
        (CI1 => CO1B) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CI0===1'b1 && CS===1'b0) 
        (CI1 => CO1B) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CI0===1'b1 && CS===1'b1) 
        (CI1 => CO1B) = (1.0, 1.0);
    ifnone
        (CI1 => CO1B) = (1.0, 1.0);

    // arc CI1 --> S
    if (A===1'b0 && B===1'b0 && CI0===1'b0) 
        (CI1 => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && CI0===1'b1) 
        (CI1 => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && CI0===1'b0) 
        (CI1 => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && CI0===1'b1) 
        (CI1 => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CI0===1'b0) 
        (CI1 => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CI0===1'b1) 
        (CI1 => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && CI0===1'b0) 
        (CI1 => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && CI0===1'b1) 
        (CI1 => S) = (1.0, 1.0);
    ifnone
        ( posedge CI1 => ( S +: CI1 ) ) = (1.0, 1.0);
        ( negedge CI1 => ( S +: CI1 ) ) = (1.0, 1.0);

    // arc CS --> S
    if (A===1'b0 && B===1'b0 && CI0===1'b0 && CI1===1'b1) 
        (CS => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && CI0===1'b1 && CI1===1'b0) 
        (CS => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && CI0===1'b0 && CI1===1'b1) 
        (CS => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && CI0===1'b1 && CI1===1'b0) 
        (CS => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CI0===1'b0 && CI1===1'b1) 
        (CS => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CI0===1'b1 && CI1===1'b0) 
        (CS => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && CI0===1'b0 && CI1===1'b1) 
        (CS => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && CI0===1'b1 && CI1===1'b0) 
        (CS => S) = (1.0, 1.0);
    ifnone
        ( posedge CS => ( S +: CS ) ) = (1.0, 1.0);
        ( negedge CS => ( S +: CS ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ADFCSOM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:02:09 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module ADFCSOM4N ( CO0B, CO1B, S, A, B, CI0, CI1, CS );
   input A, B, CI0, CI1, CS;
   output CO0B, CO1B, S;
      ADFCSOM2N_UDP5(CO0B, A, B, CI0);
      ADFCSOM2N_UDP6(CO1B, A, B, CI1);
      ADFCSOM2N_UDP7(S, A, B, CI0, CI1, CS);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO0B
    if (B===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b0) 
        (A => CO0B) = (1.0, 1.0);
    if (B===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b1) 
        (A => CO0B) = (1.0, 1.0);
    if (B===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b0) 
        (A => CO0B) = (1.0, 1.0);
    if (B===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b1) 
        (A => CO0B) = (1.0, 1.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b0) 
        (A => CO0B) = (1.0, 1.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b1) 
        (A => CO0B) = (1.0, 1.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b0) 
        (A => CO0B) = (1.0, 1.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b1) 
        (A => CO0B) = (1.0, 1.0);
    ifnone
        (A => CO0B) = (1.0, 1.0);

    // arc A --> CO1B
    if (B===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b0) 
        (A => CO1B) = (1.0, 1.0);
    if (B===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b1) 
        (A => CO1B) = (1.0, 1.0);
    if (B===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b0) 
        (A => CO1B) = (1.0, 1.0);
    if (B===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b1) 
        (A => CO1B) = (1.0, 1.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b0) 
        (A => CO1B) = (1.0, 1.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b1) 
        (A => CO1B) = (1.0, 1.0);
    if (B===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b0) 
        (A => CO1B) = (1.0, 1.0);
    if (B===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b1) 
        (A => CO1B) = (1.0, 1.0);
    ifnone
        (A => CO1B) = (1.0, 1.0);

    // arc A --> S
    if (B===1'b0 && CI0===1'b0 && CI1===1'b0 && CS===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && CI0===1'b0 && CI1===1'b0 && CS===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CI0===1'b1 && CI1===1'b1 && CS===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CI0===1'b1 && CI1===1'b1 && CS===1'b1) 
        (A => S) = (1.0, 1.0);
    ifnone
        ( posedge A => ( S +: A ) ) = (1.0, 1.0);
        ( negedge A => ( S +: A ) ) = (1.0, 1.0);

    // arc B --> CO0B
    if (A===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b0) 
        (B => CO0B) = (1.0, 1.0);
    if (A===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b1) 
        (B => CO0B) = (1.0, 1.0);
    if (A===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b0) 
        (B => CO0B) = (1.0, 1.0);
    if (A===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b1) 
        (B => CO0B) = (1.0, 1.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b0) 
        (B => CO0B) = (1.0, 1.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b1) 
        (B => CO0B) = (1.0, 1.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b0) 
        (B => CO0B) = (1.0, 1.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b1) 
        (B => CO0B) = (1.0, 1.0);
    ifnone
        (B => CO0B) = (1.0, 1.0);

    // arc B --> CO1B
    if (A===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b0) 
        (B => CO1B) = (1.0, 1.0);
    if (A===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b1) 
        (B => CO1B) = (1.0, 1.0);
    if (A===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b0) 
        (B => CO1B) = (1.0, 1.0);
    if (A===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b1) 
        (B => CO1B) = (1.0, 1.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b0) 
        (B => CO1B) = (1.0, 1.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b1) 
        (B => CO1B) = (1.0, 1.0);
    if (A===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b0) 
        (B => CO1B) = (1.0, 1.0);
    if (A===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b1) 
        (B => CO1B) = (1.0, 1.0);
    ifnone
        (B => CO1B) = (1.0, 1.0);

    // arc B --> S
    if (A===1'b0 && CI0===1'b0 && CI1===1'b0 && CS===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && CI0===1'b0 && CI1===1'b0 && CS===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CI0===1'b1 && CI1===1'b1 && CS===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CI0===1'b1 && CI1===1'b1 && CS===1'b1) 
        (B => S) = (1.0, 1.0);
    ifnone
        ( posedge B => ( S +: B ) ) = (1.0, 1.0);
        ( negedge B => ( S +: B ) ) = (1.0, 1.0);

    // arc CI0 --> CO0B
    if (A===1'b0 && B===1'b1 && CI1===1'b0 && CS===1'b0) 
        (CI0 => CO0B) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && CI1===1'b0 && CS===1'b1) 
        (CI0 => CO0B) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && CI1===1'b1 && CS===1'b0) 
        (CI0 => CO0B) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && CI1===1'b1 && CS===1'b1) 
        (CI0 => CO0B) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CI1===1'b0 && CS===1'b0) 
        (CI0 => CO0B) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CI1===1'b0 && CS===1'b1) 
        (CI0 => CO0B) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CI1===1'b1 && CS===1'b0) 
        (CI0 => CO0B) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CI1===1'b1 && CS===1'b1) 
        (CI0 => CO0B) = (1.0, 1.0);
    ifnone
        (CI0 => CO0B) = (1.0, 1.0);

    // arc CI0 --> S
    if (A===1'b0 && B===1'b0 && CI1===1'b0) 
        (CI0 => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && CI1===1'b1) 
        (CI0 => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && CI1===1'b0) 
        (CI0 => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && CI1===1'b1) 
        (CI0 => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CI1===1'b0) 
        (CI0 => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CI1===1'b1) 
        (CI0 => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && CI1===1'b0) 
        (CI0 => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && CI1===1'b1) 
        (CI0 => S) = (1.0, 1.0);
    ifnone
        ( posedge CI0 => ( S +: CI0 ) ) = (1.0, 1.0);
        ( negedge CI0 => ( S +: CI0 ) ) = (1.0, 1.0);

    // arc CI1 --> CO1B
    if (A===1'b0 && B===1'b1 && CI0===1'b0 && CS===1'b0) 
        (CI1 => CO1B) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && CI0===1'b0 && CS===1'b1) 
        (CI1 => CO1B) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && CI0===1'b1 && CS===1'b0) 
        (CI1 => CO1B) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && CI0===1'b1 && CS===1'b1) 
        (CI1 => CO1B) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CI0===1'b0 && CS===1'b0) 
        (CI1 => CO1B) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CI0===1'b0 && CS===1'b1) 
        (CI1 => CO1B) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CI0===1'b1 && CS===1'b0) 
        (CI1 => CO1B) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CI0===1'b1 && CS===1'b1) 
        (CI1 => CO1B) = (1.0, 1.0);
    ifnone
        (CI1 => CO1B) = (1.0, 1.0);

    // arc CI1 --> S
    if (A===1'b0 && B===1'b0 && CI0===1'b0) 
        (CI1 => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && CI0===1'b1) 
        (CI1 => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && CI0===1'b0) 
        (CI1 => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && CI0===1'b1) 
        (CI1 => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CI0===1'b0) 
        (CI1 => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CI0===1'b1) 
        (CI1 => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && CI0===1'b0) 
        (CI1 => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && CI0===1'b1) 
        (CI1 => S) = (1.0, 1.0);
    ifnone
        ( posedge CI1 => ( S +: CI1 ) ) = (1.0, 1.0);
        ( negedge CI1 => ( S +: CI1 ) ) = (1.0, 1.0);

    // arc CS --> S
    if (A===1'b0 && B===1'b0 && CI0===1'b0 && CI1===1'b1) 
        (CS => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && CI0===1'b1 && CI1===1'b0) 
        (CS => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && CI0===1'b0 && CI1===1'b1) 
        (CS => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && CI0===1'b1 && CI1===1'b0) 
        (CS => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CI0===1'b0 && CI1===1'b1) 
        (CS => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && CI0===1'b1 && CI1===1'b0) 
        (CS => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && CI0===1'b0 && CI1===1'b1) 
        (CS => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && CI0===1'b1 && CI1===1'b0) 
        (CS => S) = (1.0, 1.0);
    ifnone
        ( posedge CS => ( S +: CS ) ) = (1.0, 1.0);
        ( negedge CS => ( S +: CS ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ADFCSOM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:02:43 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module ADFM0N ( CO, S, A, B, CI );
   input A, B, CI;
   output CO, S;
      ADFM0N_UDP3(CO, A, B, CI);
      ADFM0N_UDP4(S, A, B, CI);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO
    if (B===1'b0 && CI===1'b1) 
        (A => CO) = (1.0, 1.0);
    if (B===1'b1 && CI===1'b0) 
        (A => CO) = (1.0, 1.0);
    ifnone
        (A => CO) = (1.0, 1.0);

    // arc A --> S
    if (B===1'b0 && CI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && CI===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CI===1'b1) 
        (A => S) = (1.0, 1.0);
    ifnone
        ( posedge A => ( S +: A ) ) = (1.0, 1.0);
        ( negedge A => ( S +: A ) ) = (1.0, 1.0);

    // arc B --> CO
    if (A===1'b0 && CI===1'b1) 
        (B => CO) = (1.0, 1.0);
    if (A===1'b1 && CI===1'b0) 
        (B => CO) = (1.0, 1.0);
    ifnone
        (B => CO) = (1.0, 1.0);

    // arc B --> S
    if (A===1'b0 && CI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && CI===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CI===1'b1) 
        (B => S) = (1.0, 1.0);
    ifnone
        ( posedge B => ( S +: B ) ) = (1.0, 1.0);
        ( negedge B => ( S +: B ) ) = (1.0, 1.0);

    // arc CI --> CO
    if (A===1'b0 && B===1'b1) 
        (CI => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0) 
        (CI => CO) = (1.0, 1.0);
    ifnone
        (CI => CO) = (1.0, 1.0);

    // arc CI --> S
    if (A===1'b0 && B===1'b0) 
        (CI => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1) 
        (CI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0) 
        (CI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1) 
        (CI => S) = (1.0, 1.0);
    ifnone
        ( posedge CI => ( S +: CI ) ) = (1.0, 1.0);
        ( negedge CI => ( S +: CI ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ADFM0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:03:42 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module ADFM1N ( CO, S, A, B, CI );
   input A, B, CI;
   output CO, S;
      ADFM0N_UDP3(CO, A, B, CI);
      ADFM0N_UDP4(S, A, B, CI);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO
    if (B===1'b0 && CI===1'b1) 
        (A => CO) = (1.0, 1.0);
    if (B===1'b1 && CI===1'b0) 
        (A => CO) = (1.0, 1.0);
    ifnone
        (A => CO) = (1.0, 1.0);

    // arc A --> S
    if (B===1'b0 && CI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && CI===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CI===1'b1) 
        (A => S) = (1.0, 1.0);
    ifnone
        ( posedge A => ( S +: A ) ) = (1.0, 1.0);
        ( negedge A => ( S +: A ) ) = (1.0, 1.0);

    // arc B --> CO
    if (A===1'b0 && CI===1'b1) 
        (B => CO) = (1.0, 1.0);
    if (A===1'b1 && CI===1'b0) 
        (B => CO) = (1.0, 1.0);
    ifnone
        (B => CO) = (1.0, 1.0);

    // arc B --> S
    if (A===1'b0 && CI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && CI===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CI===1'b1) 
        (B => S) = (1.0, 1.0);
    ifnone
        ( posedge B => ( S +: B ) ) = (1.0, 1.0);
        ( negedge B => ( S +: B ) ) = (1.0, 1.0);

    // arc CI --> CO
    if (A===1'b0 && B===1'b1) 
        (CI => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0) 
        (CI => CO) = (1.0, 1.0);
    ifnone
        (CI => CO) = (1.0, 1.0);

    // arc CI --> S
    if (A===1'b0 && B===1'b0) 
        (CI => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1) 
        (CI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0) 
        (CI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1) 
        (CI => S) = (1.0, 1.0);
    ifnone
        ( posedge CI => ( S +: CI ) ) = (1.0, 1.0);
        ( negedge CI => ( S +: CI ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ADFM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:07:31 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module ADFM2N ( CO, S, A, B, CI );
   input A, B, CI;
   output CO, S;
      ADFM0N_UDP3(CO, A, B, CI);
      ADFM0N_UDP4(S, A, B, CI);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO
    if (B===1'b0 && CI===1'b1) 
        (A => CO) = (1.0, 1.0);
    if (B===1'b1 && CI===1'b0) 
        (A => CO) = (1.0, 1.0);
    ifnone
        (A => CO) = (1.0, 1.0);

    // arc A --> S
    if (B===1'b0 && CI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && CI===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CI===1'b1) 
        (A => S) = (1.0, 1.0);
    ifnone
        ( posedge A => ( S +: A ) ) = (1.0, 1.0);
        ( negedge A => ( S +: A ) ) = (1.0, 1.0);

    // arc B --> CO
    if (A===1'b0 && CI===1'b1) 
        (B => CO) = (1.0, 1.0);
    if (A===1'b1 && CI===1'b0) 
        (B => CO) = (1.0, 1.0);
    ifnone
        (B => CO) = (1.0, 1.0);

    // arc B --> S
    if (A===1'b0 && CI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && CI===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CI===1'b1) 
        (B => S) = (1.0, 1.0);
    ifnone
        ( posedge B => ( S +: B ) ) = (1.0, 1.0);
        ( negedge B => ( S +: B ) ) = (1.0, 1.0);

    // arc CI --> CO
    if (A===1'b0 && B===1'b1) 
        (CI => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0) 
        (CI => CO) = (1.0, 1.0);
    ifnone
        (CI => CO) = (1.0, 1.0);

    // arc CI --> S
    if (A===1'b0 && B===1'b0) 
        (CI => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1) 
        (CI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0) 
        (CI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1) 
        (CI => S) = (1.0, 1.0);
    ifnone
        ( posedge CI => ( S +: CI ) ) = (1.0, 1.0);
        ( negedge CI => ( S +: CI ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ADFM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:08:57 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module ADFM4N ( CO, S, A, B, CI );
   input A, B, CI;
   output CO, S;
      ADFM0N_UDP3(CO, A, B, CI);
      ADFM0N_UDP4(S, A, B, CI);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO
    if (B===1'b0 && CI===1'b1) 
        (A => CO) = (1.0, 1.0);
    if (B===1'b1 && CI===1'b0) 
        (A => CO) = (1.0, 1.0);
    ifnone
        (A => CO) = (1.0, 1.0);

    // arc A --> S
    if (B===1'b0 && CI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && CI===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CI===1'b1) 
        (A => S) = (1.0, 1.0);
    ifnone
        ( posedge A => ( S +: A ) ) = (1.0, 1.0);
        ( negedge A => ( S +: A ) ) = (1.0, 1.0);

    // arc B --> CO
    if (A===1'b0 && CI===1'b1) 
        (B => CO) = (1.0, 1.0);
    if (A===1'b1 && CI===1'b0) 
        (B => CO) = (1.0, 1.0);
    ifnone
        (B => CO) = (1.0, 1.0);

    // arc B --> S
    if (A===1'b0 && CI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && CI===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CI===1'b1) 
        (B => S) = (1.0, 1.0);
    ifnone
        ( posedge B => ( S +: B ) ) = (1.0, 1.0);
        ( negedge B => ( S +: B ) ) = (1.0, 1.0);

    // arc CI --> CO
    if (A===1'b0 && B===1'b1) 
        (CI => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0) 
        (CI => CO) = (1.0, 1.0);
    ifnone
        (CI => CO) = (1.0, 1.0);

    // arc CI --> S
    if (A===1'b0 && B===1'b0) 
        (CI => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1) 
        (CI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0) 
        (CI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1) 
        (CI => S) = (1.0, 1.0);
    ifnone
        ( posedge CI => ( S +: CI ) ) = (1.0, 1.0);
        ( negedge CI => ( S +: CI ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ADFM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:05:13 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module ADFOM2N ( COB, S, A, B, CI );
   input A, B, CI;
   output COB, S;
      ADFOM2N_UDP3(COB, A, B, CI);
      ADFOM2N_UDP4(S, A, B, CI);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> COB
    if (B===1'b0 && CI===1'b1) 
        (A => COB) = (1.0, 1.0);
    if (B===1'b1 && CI===1'b0) 
        (A => COB) = (1.0, 1.0);
    ifnone
        (A => COB) = (1.0, 1.0);

    // arc A --> S
    if (B===1'b0 && CI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && CI===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CI===1'b1) 
        (A => S) = (1.0, 1.0);
    ifnone
        ( posedge A => ( S +: A ) ) = (1.0, 1.0);
        ( negedge A => ( S +: A ) ) = (1.0, 1.0);

    // arc B --> COB
    if (A===1'b0 && CI===1'b1) 
        (B => COB) = (1.0, 1.0);
    if (A===1'b1 && CI===1'b0) 
        (B => COB) = (1.0, 1.0);
    ifnone
        (B => COB) = (1.0, 1.0);

    // arc B --> S
    if (A===1'b0 && CI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && CI===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CI===1'b1) 
        (B => S) = (1.0, 1.0);
    ifnone
        ( posedge B => ( S +: B ) ) = (1.0, 1.0);
        ( negedge B => ( S +: B ) ) = (1.0, 1.0);

    // arc CI --> COB
    if (A===1'b0 && B===1'b1) 
        (CI => COB) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0) 
        (CI => COB) = (1.0, 1.0);
    ifnone
        (CI => COB) = (1.0, 1.0);

    // arc CI --> S
    if (A===1'b0 && B===1'b0) 
        (CI => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1) 
        (CI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0) 
        (CI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1) 
        (CI => S) = (1.0, 1.0);
    ifnone
        ( posedge CI => ( S +: CI ) ) = (1.0, 1.0);
        ( negedge CI => ( S +: CI ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ADFOM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:08:33 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module ADFOM4N ( COB, S, A, B, CI );
   input A, B, CI;
   output COB, S;
      ADFOM2N_UDP3(COB, A, B, CI);
      ADFOM2N_UDP4(S, A, B, CI);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> COB
    if (B===1'b0 && CI===1'b1) 
        (A => COB) = (1.0, 1.0);
    if (B===1'b1 && CI===1'b0) 
        (A => COB) = (1.0, 1.0);
    ifnone
        (A => COB) = (1.0, 1.0);

    // arc A --> S
    if (B===1'b0 && CI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && CI===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CI===1'b1) 
        (A => S) = (1.0, 1.0);
    ifnone
        ( posedge A => ( S +: A ) ) = (1.0, 1.0);
        ( negedge A => ( S +: A ) ) = (1.0, 1.0);

    // arc B --> COB
    if (A===1'b0 && CI===1'b1) 
        (B => COB) = (1.0, 1.0);
    if (A===1'b1 && CI===1'b0) 
        (B => COB) = (1.0, 1.0);
    ifnone
        (B => COB) = (1.0, 1.0);

    // arc B --> S
    if (A===1'b0 && CI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && CI===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CI===1'b1) 
        (B => S) = (1.0, 1.0);
    ifnone
        ( posedge B => ( S +: B ) ) = (1.0, 1.0);
        ( negedge B => ( S +: B ) ) = (1.0, 1.0);

    // arc CI --> COB
    if (A===1'b0 && B===1'b1) 
        (CI => COB) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0) 
        (CI => COB) = (1.0, 1.0);
    ifnone
        (CI => COB) = (1.0, 1.0);

    // arc CI --> S
    if (A===1'b0 && B===1'b0) 
        (CI => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1) 
        (CI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0) 
        (CI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1) 
        (CI => S) = (1.0, 1.0);
    ifnone
        ( posedge CI => ( S +: CI ) ) = (1.0, 1.0);
        ( negedge CI => ( S +: CI ) ) = (1.0, 1.0);



  endspecify
  `endif // functional //
endmodule     // ADFOM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:03:01 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADHCM2N(A, NCI, CO, S);
  input A, NCI;
  output CO, S;

    not SMC_I0(NCI_bar, NCI);
    and SMC_I1(CO, A, NCI_bar);

    xnor SMC_I2(S, A, NCI);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO
    (A => CO) = (1.0, 1.0);

    // arc A --> S
     if ( A===1'b1 )
    ( posedge A => ( S +: A ) ) = (1.0, 1.0);
     if ( A===1'b0 )
    ( negedge A => ( S +: A ) ) = (1.0, 1.0);

    // arc NCI --> CO
    (NCI => CO) = (1.0, 1.0);

    // arc NCI --> S
     if ( NCI===1'b1 )
    ( posedge NCI => ( S +: NCI ) ) = (1.0, 1.0);
     if ( NCI===1'b0 )
    ( negedge NCI => ( S +: NCI ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ADHCM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:05:59 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADHCM4N(A, NCI, CO, S);
  input A, NCI;
  output CO, S;

    not SMC_I0(NCI_bar, NCI);
    and SMC_I1(CO, A, NCI_bar);

    xnor SMC_I2(S, A, NCI);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO
    (A => CO) = (1.0, 1.0);

    // arc A --> S
     if ( A===1'b1 )
    ( posedge A => ( S +: A ) ) = (1.0, 1.0);
     if ( A===1'b0 )
    ( negedge A => ( S +: A ) ) = (1.0, 1.0);

    // arc NCI --> CO
    (NCI => CO) = (1.0, 1.0);

    // arc NCI --> S
     if ( NCI===1'b1 )
    ( posedge NCI => ( S +: NCI ) ) = (1.0, 1.0);
     if ( NCI===1'b0 )
    ( negedge NCI => ( S +: NCI ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ADHCM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:10:10 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADHCSCM2N(A, CS, NCI, CO, S);
  input A, CS, NCI;
  output CO, S;

    not SMC_I0(NCI_bar, NCI);
    and SMC_I1(CO, A, NCI_bar);

    not SMC_I2(A_bar, A);
    and SMC_I3(OUT0, A_bar, CS, NCI_bar);
    not SMC_I4(CS_bar, CS);
    and SMC_I5(OUT1, A, CS_bar);
    and SMC_I6(OUT2, A, NCI);
    or SMC_I7(S, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO
    if (CS===1'b0) 
        (A => CO) = (1.0, 1.0);
    if (CS===1'b1) 
        (A => CO) = (1.0, 1.0);
    ifnone
        (A => CO) = (1.0, 1.0);

    // arc A --> S
    if (CS===1'b0 && NCI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (CS===1'b0 && NCI===1'b1) 
        (A => S) = (1.0, 1.0);
    if (CS===1'b1 && NCI===1'b1) 
        (A => S) = (1.0, 1.0);
    ifnone
        ( posedge A => ( S +: A ) ) = (1.0, 1.0);
        ( negedge A => ( S +: A ) ) = (1.0, 1.0);

    // arc CS --> S
     if ( CS===1'b1 )
    ( posedge CS => ( S +: CS ) ) = (1.0, 1.0);
     if ( CS===1'b0 )
    ( negedge CS => ( S +: CS ) ) = (1.0, 1.0);

    // arc NCI --> CO
    if (CS===1'b0) 
        (NCI => CO) = (1.0, 1.0);
    if (CS===1'b1) 
        (NCI => CO) = (1.0, 1.0);
    ifnone
        (NCI => CO) = (1.0, 1.0);

    // arc NCI --> S
     if ( NCI===1'b1 )
    ( posedge NCI => ( S +: NCI ) ) = (1.0, 1.0);
     if ( NCI===1'b0 )
    ( negedge NCI => ( S +: NCI ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ADHCSCM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:08:09 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADHCSCM4N(A, CS, NCI, CO, S);
  input A, CS, NCI;
  output CO, S;

    not SMC_I0(NCI_bar, NCI);
    and SMC_I1(CO, A, NCI_bar);

    not SMC_I2(A_bar, A);
    and SMC_I3(OUT0, A_bar, CS, NCI_bar);
    not SMC_I4(CS_bar, CS);
    and SMC_I5(OUT1, A, CS_bar);
    and SMC_I6(OUT2, A, NCI);
    or SMC_I7(S, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO
    if (CS===1'b0) 
        (A => CO) = (1.0, 1.0);
    if (CS===1'b1) 
        (A => CO) = (1.0, 1.0);
    ifnone
        (A => CO) = (1.0, 1.0);

    // arc A --> S
    if (CS===1'b0 && NCI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (CS===1'b0 && NCI===1'b1) 
        (A => S) = (1.0, 1.0);
    if (CS===1'b1 && NCI===1'b1) 
        (A => S) = (1.0, 1.0);
    ifnone
        ( posedge A => ( S +: A ) ) = (1.0, 1.0);
        ( negedge A => ( S +: A ) ) = (1.0, 1.0);

    // arc CS --> S
     if ( CS===1'b1 )
    ( posedge CS => ( S +: CS ) ) = (1.0, 1.0);
     if ( CS===1'b0 )
    ( negedge CS => ( S +: CS ) ) = (1.0, 1.0);

    // arc NCI --> CO
    if (CS===1'b0) 
        (NCI => CO) = (1.0, 1.0);
    if (CS===1'b1) 
        (NCI => CO) = (1.0, 1.0);
    ifnone
        (NCI => CO) = (1.0, 1.0);

    // arc NCI --> S
     if ( NCI===1'b1 )
    ( posedge NCI => ( S +: NCI ) ) = (1.0, 1.0);
     if ( NCI===1'b0 )
    ( negedge NCI => ( S +: NCI ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ADHCSCM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:03:05 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADHCSOM2N(A, CI, CS, COB, S);
  input A, CI, CS;
  output COB, S;

    nand SMC_I0(COB, A, CI);

    not SMC_I1(CS_bar, CS);
    and SMC_I2(OUT0, A, CS_bar);
    not SMC_I3(CI_bar, CI);
    and SMC_I4(OUT1, A, CI_bar);
    not SMC_I5(A_bar, A);
    and SMC_I6(OUT2, A_bar, CI, CS);
    or SMC_I7(S, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> COB
    if (CS===1'b0) 
        (A => COB) = (1.0, 1.0);
    if (CS===1'b1) 
        (A => COB) = (1.0, 1.0);
    ifnone
        (A => COB) = (1.0, 1.0);

    // arc A --> S
    if (CI===1'b0 && CS===1'b0) 
        (A => S) = (1.0, 1.0);
    if (CI===1'b0 && CS===1'b1) 
        (A => S) = (1.0, 1.0);
    if (CI===1'b1 && CS===1'b0) 
        (A => S) = (1.0, 1.0);
    ifnone
        ( posedge A => ( S +: A ) ) = (1.0, 1.0);
        ( negedge A => ( S +: A ) ) = (1.0, 1.0);

    // arc CI --> COB
    if (CS===1'b0) 
        (CI => COB) = (1.0, 1.0);
    if (CS===1'b1) 
        (CI => COB) = (1.0, 1.0);
    ifnone
        (CI => COB) = (1.0, 1.0);

    // arc CI --> S
     if ( CI===1'b1 )
    ( posedge CI => ( S +: CI ) ) = (1.0, 1.0);
     if ( CI===1'b0 )
    ( negedge CI => ( S +: CI ) ) = (1.0, 1.0);

    // arc CS --> S
     if ( CS===1'b1 )
    ( posedge CS => ( S +: CS ) ) = (1.0, 1.0);
     if ( CS===1'b0 )
    ( negedge CS => ( S +: CS ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ADHCSOM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:06:10 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADHCSOM4N(A, CI, CS, COB, S);
  input A, CI, CS;
  output COB, S;

    nand SMC_I0(COB, A, CI);

    not SMC_I1(CS_bar, CS);
    and SMC_I2(OUT0, A, CS_bar);
    not SMC_I3(CI_bar, CI);
    and SMC_I4(OUT1, A, CI_bar);
    not SMC_I5(A_bar, A);
    and SMC_I6(OUT2, A_bar, CI, CS);
    or SMC_I7(S, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> COB
    if (CS===1'b0) 
        (A => COB) = (1.0, 1.0);
    if (CS===1'b1) 
        (A => COB) = (1.0, 1.0);
    ifnone
        (A => COB) = (1.0, 1.0);

    // arc A --> S
    if (CI===1'b0 && CS===1'b0) 
        (A => S) = (1.0, 1.0);
    if (CI===1'b0 && CS===1'b1) 
        (A => S) = (1.0, 1.0);
    if (CI===1'b1 && CS===1'b0) 
        (A => S) = (1.0, 1.0);
    ifnone
        ( posedge A => ( S +: A ) ) = (1.0, 1.0);
        ( negedge A => ( S +: A ) ) = (1.0, 1.0);

    // arc CI --> COB
    if (CS===1'b0) 
        (CI => COB) = (1.0, 1.0);
    if (CS===1'b1) 
        (CI => COB) = (1.0, 1.0);
    ifnone
        (CI => COB) = (1.0, 1.0);

    // arc CI --> S
     if ( CI===1'b1 )
    ( posedge CI => ( S +: CI ) ) = (1.0, 1.0);
     if ( CI===1'b0 )
    ( negedge CI => ( S +: CI ) ) = (1.0, 1.0);

    // arc CS --> S
     if ( CS===1'b1 )
    ( posedge CS => ( S +: CS ) ) = (1.0, 1.0);
     if ( CS===1'b0 )
    ( negedge CS => ( S +: CS ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ADHCSOM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:03:51 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADHM0N(A, B, CO, S);
  input A, B;
  output CO, S;

    and SMC_I0(CO, A, B);

    xor SMC_I1(S, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO
    (A => CO) = (1.0, 1.0);

    // arc A --> S
     if ( A===1'b1 )
    ( posedge A => ( S +: A ) ) = (1.0, 1.0);
     if ( A===1'b0 )
    ( negedge A => ( S +: A ) ) = (1.0, 1.0);

    // arc B --> CO
    (B => CO) = (1.0, 1.0);

    // arc B --> S
     if ( B===1'b1 )
    ( posedge B => ( S +: B ) ) = (1.0, 1.0);
     if ( B===1'b0 )
    ( negedge B => ( S +: B ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ADHM0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:08:41 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADHM1N(A, B, CO, S);
  input A, B;
  output CO, S;

    and SMC_I0(CO, A, B);

    xor SMC_I1(S, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO
    (A => CO) = (1.0, 1.0);

    // arc A --> S
     if ( A===1'b1 )
    ( posedge A => ( S +: A ) ) = (1.0, 1.0);
     if ( A===1'b0 )
    ( negedge A => ( S +: A ) ) = (1.0, 1.0);

    // arc B --> CO
    (B => CO) = (1.0, 1.0);

    // arc B --> S
     if ( B===1'b1 )
    ( posedge B => ( S +: B ) ) = (1.0, 1.0);
     if ( B===1'b0 )
    ( negedge B => ( S +: B ) ) = (1.0, 1.0);



  endspecify
  `endif // functional //
endmodule     // ADHM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:05:37 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADHM2N(A, B, CO, S);
  input A, B;
  output CO, S;

    and SMC_I0(CO, A, B);

    xor SMC_I1(S, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO
    (A => CO) = (1.0, 1.0);

    // arc A --> S
     if ( A===1'b1 )
    ( posedge A => ( S +: A ) ) = (1.0, 1.0);
     if ( A===1'b0 )
    ( negedge A => ( S +: A ) ) = (1.0, 1.0);

    // arc B --> CO
    (B => CO) = (1.0, 1.0);

    // arc B --> S
     if ( B===1'b1 )
    ( posedge B => ( S +: B ) ) = (1.0, 1.0);
     if ( B===1'b0 )
    ( negedge B => ( S +: B ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ADHM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:10:20 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADHM4N(A, B, CO, S);
  input A, B;
  output CO, S;

    and SMC_I0(CO, A, B);

    xor SMC_I1(S, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO
    (A => CO) = (1.0, 1.0);

    // arc A --> S
     if ( A===1'b1 )
    ( posedge A => ( S +: A ) ) = (1.0, 1.0);
     if ( A===1'b0 )
    ( negedge A => ( S +: A ) ) = (1.0, 1.0);

    // arc B --> CO
    (B => CO) = (1.0, 1.0);

    // arc B --> S
     if ( B===1'b1 )
    ( posedge B => ( S +: B ) ) = (1.0, 1.0);
     if ( B===1'b0 )
    ( negedge B => ( S +: B ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ADHM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:07:52 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADHOM2N(A, CI, COB, S);
  input A, CI;
  output COB, S;

    nand SMC_I0(COB, A, CI);

    xor SMC_I1(S, A, CI);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> COB
    (A => COB) = (1.0, 1.0);

    // arc A --> S
     if ( A===1'b1 )
    ( posedge A => ( S +: A ) ) = (1.0, 1.0);
     if ( A===1'b0 )
    ( negedge A => ( S +: A ) ) = (1.0, 1.0);

    // arc CI --> COB
    (CI => COB) = (1.0, 1.0);

    // arc CI --> S
     if ( CI===1'b1 )
    ( posedge CI => ( S +: CI ) ) = (1.0, 1.0);
     if ( CI===1'b0 )
    ( negedge CI => ( S +: CI ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ADHOM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:09:15 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADHOM4N(A, CI, COB, S);
  input A, CI;
  output COB, S;

    nand SMC_I0(COB, A, CI);

    xor SMC_I1(S, A, CI);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> COB
    (A => COB) = (1.0, 1.0);

    // arc A --> S
     if ( A===1'b1 )
    ( posedge A => ( S +: A ) ) = (1.0, 1.0);
     if ( A===1'b0 )
    ( negedge A => ( S +: A ) ) = (1.0, 1.0);

    // arc CI --> COB
    (CI => COB) = (1.0, 1.0);

    // arc CI --> S
     if ( CI===1'b1 )
    ( posedge CI => ( S +: CI ) ) = (1.0, 1.0);
     if ( CI===1'b0 )
    ( negedge CI => ( S +: CI ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ADHOM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:08:21 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AN2M0N(A, B, Z);
  input A, B;
  output Z;

    and SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AN2M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:03:59 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AN2M1N(A, B, Z);
  input A, B;
  output Z;

    and SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AN2M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:06:31 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AN2M2N(A, B, Z);
  input A, B;
  output Z;

    and SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AN2M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:08:05 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AN2M4N(A, B, Z);
  input A, B;
  output Z;

    and SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AN2M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:05:38 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AN2M6N(A, B, Z);
  input A, B;
  output Z;

    and SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AN2M6N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:07:01 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AN2M8N(A, B, Z);
  input A, B;
  output Z;

    and SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AN2M8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:06:16 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module AN3M0N ( Z, A, B, C );
   input A, B, C;
   output Z;
      AN3M0N_UDP3(Z, A, B, C);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AN3M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:08:48 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module AN3M1N ( Z, A, B, C );
   input A, B, C;
   output Z;
      AN3M0N_UDP3(Z, A, B, C);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AN3M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:07:16 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module AN3M2N ( Z, A, B, C );
   input A, B, C;
   output Z;
      AN3M0N_UDP3(Z, A, B, C);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AN3M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:08:20 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module AN3M4N ( Z, A, B, C );
   input A, B, C;
   output Z;
      AN3M0N_UDP3(Z, A, B, C);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AN3M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:05:53 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module AN3M6N ( Z, A, B, C );
   input A, B, C;
   output Z;
      AN3M0N_UDP3(Z, A, B, C);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AN3M6N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:04:14 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module AN3M8N ( Z, A, B, C );
   input A, B, C;
   output Z;
      AN3M0N_UDP3(Z, A, B, C);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AN3M8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:06:46 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module AN4M0N ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;
      AN4M0N_UDP4(Z, A, B, C, D);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc D --> Z
    (D => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AN4M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:01:30 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module AN4M1N ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;
      AN4M0N_UDP4(Z, A, B, C, D);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc D --> Z
    (D => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AN4M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:03:54 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module AN4M2N ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;
      AN4M0N_UDP4(Z, A, B, C, D);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc D --> Z
    (D => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AN4M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:07:31 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module AN4M4N ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;
      AN4M0N_UDP4(Z, A, B, C, D);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc D --> Z
    (D => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AN4M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:08:35 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module AN4M6N ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;
      AN4M0N_UDP4(Z, A, B, C, D);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc D --> Z
    (D => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AN4M6N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:06:08 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module AN4M8N ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;
      AN4M0N_UDP4(Z, A, B, C, D);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc D --> Z
    (D => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AN4M8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:04:09 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO21M0N(A1, A2, B, Z);
  input A1, A2, B;
  output Z;

    and SMC_I0(OUT0, A1, A2);
    buf SMC_I1(OUT1, B);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AO21M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:06:23 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO21M1N(A1, A2, B, Z);
  input A1, A2, B;
  output Z;

    and SMC_I0(OUT0, A1, A2);
    buf SMC_I1(OUT1, B);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AO21M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:01:42 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO21M2N(A1, A2, B, Z);
  input A1, A2, B;
  output Z;

    and SMC_I0(OUT0, A1, A2);
    buf SMC_I1(OUT1, B);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AO21M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:01:45 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO21M4N(A1, A2, B, Z);
  input A1, A2, B;
  output Z;

    and SMC_I0(OUT0, A1, A2);
    buf SMC_I1(OUT1, B);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AO21M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:01:45 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module AO22B10M0N ( Z, A1, B1, B2, NA2 );
   input A1, B1, B2, NA2;
   output Z;
      AO22B10M0N_UDP4(Z, A1, B1, B2, NA2);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);

    // arc NA2 --> Z
    (NA2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AO22B10M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:03:17 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module AO22B10M1N ( Z, A1, B1, B2, NA2 );
   input A1, B1, B2, NA2;
   output Z;
      AO22B10M0N_UDP4(Z, A1, B1, B2, NA2);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);

    // arc NA2 --> Z
    (NA2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AO22B10M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:07:46 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module AO22B10M2N ( Z, A1, B1, B2, NA2 );
   input A1, B1, B2, NA2;
   output Z;
      AO22B10M0N_UDP4(Z, A1, B1, B2, NA2);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);

    // arc NA2 --> Z
    (NA2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AO22B10M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:08:24 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module AO22B10M4N ( Z, A1, B1, B2, NA2 );
   input A1, B1, B2, NA2;
   output Z;
      AO22B10M0N_UDP4(Z, A1, B1, B2, NA2);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);

    // arc NA2 --> Z
    (NA2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AO22B10M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:04:24 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module AO22B11M0N ( Z, A1, B1, NA2, NB2 );
   input A1, B1, NA2, NB2;
   output Z;
      AO22B11M0N_UDP4(Z, A1, B1, NA2, NB2);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc NA2 --> Z
    (NA2 => Z) = (1.0, 1.0);

    // arc NB2 --> Z
    (NB2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AO22B11M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:06:38 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module AO22B11M1N ( Z, A1, B1, NA2, NB2 );
   input A1, B1, NA2, NB2;
   output Z;
      AO22B11M0N_UDP4(Z, A1, B1, NA2, NB2);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc NA2 --> Z
    (NA2 => Z) = (1.0, 1.0);

    // arc NB2 --> Z
    (NB2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AO22B11M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:01:59 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module AO22B11M2N ( Z, A1, B1, NA2, NB2 );
   input A1, B1, NA2, NB2;
   output Z;
      AO22B11M0N_UDP4(Z, A1, B1, NA2, NB2);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc NA2 --> Z
    (NA2 => Z) = (1.0, 1.0);

    // arc NB2 --> Z
    (NB2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AO22B11M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:01:57 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module AO22B11M4N ( Z, A1, B1, NA2, NB2 );
   input A1, B1, NA2, NB2;
   output Z;
      AO22B11M0N_UDP4(Z, A1, B1, NA2, NB2);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc NA2 --> Z
    (NA2 => Z) = (1.0, 1.0);

    // arc NB2 --> Z
    (NB2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AO22B11M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:02:00 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module AO22M0N ( Z, A1, A2, B1, B2 );
   input A1, A2, B1, B2;
   output Z;
      AO22M0N_UDP4(Z, A1, A2, B1, B2);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AO22M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:09:05 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module AO22M1N ( Z, A1, A2, B1, B2 );
   input A1, A2, B1, B2;
   output Z;
      AO22M0N_UDP4(Z, A1, A2, B1, B2);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AO22M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:06:21 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module AO22M2N ( Z, A1, A2, B1, B2 );
   input A1, A2, B1, B2;
   output Z;
      AO22M0N_UDP4(Z, A1, A2, B1, B2);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AO22M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:09:23 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module AO22M4N ( Z, A1, A2, B1, B2 );
   input A1, A2, B1, B2;
   output Z;
      AO22M0N_UDP4(Z, A1, A2, B1, B2);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AO22M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:08:56 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI211M0N ( Z, A1, A2, B, C );
   input A1, A2, B, C;
   output Z;
      AOI211M0N_UDP4(Z, A1, A2, B, C);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI211M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:05:49 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI211M1N ( Z, A1, A2, B, C );
   input A1, A2, B, C;
   output Z;
      AOI211M0N_UDP4(Z, A1, A2, B, C);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI211M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:08:06 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI211M2N ( Z, A1, A2, B, C );
   input A1, A2, B, C;
   output Z;
      AOI211M0N_UDP4(Z, A1, A2, B, C);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI211M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:04:12 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI211M4N ( Z, A1, A2, B, C );
   input A1, A2, B, C;
   output Z;
      AOI211M0N_UDP4(Z, A1, A2, B, C);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI211M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:02:16 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21B01M0N(A1, A2, NB, Z);
  input A1, A2, NB;
  output Z;

    not SMC_I0(A1_bar, A1);
    and SMC_I1(OUT0, A1_bar, NB);
    not SMC_I2(A2_bar, A2);
    and SMC_I3(OUT1, A2_bar, NB);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc NB --> Z
    (NB => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI21B01M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:09:21 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21B01M1N(A1, A2, NB, Z);
  input A1, A2, NB;
  output Z;

    not SMC_I0(A1_bar, A1);
    and SMC_I1(OUT0, A1_bar, NB);
    not SMC_I2(A2_bar, A2);
    and SMC_I3(OUT1, A2_bar, NB);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc NB --> Z
    (NB => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI21B01M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:02:14 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21B01M2N(A1, A2, NB, Z);
  input A1, A2, NB;
  output Z;

    not SMC_I0(A1_bar, A1);
    and SMC_I1(OUT0, A1_bar, NB);
    not SMC_I2(A2_bar, A2);
    and SMC_I3(OUT1, A2_bar, NB);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc NB --> Z
    (NB => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI21B01M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:02:16 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21B01M4N(A1, A2, NB, Z);
  input A1, A2, NB;
  output Z;

    not SMC_I0(A1_bar, A1);
    and SMC_I1(OUT0, A1_bar, NB);
    not SMC_I2(A2_bar, A2);
    and SMC_I3(OUT1, A2_bar, NB);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc NB --> Z
    (NB => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI21B01M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:04:41 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21B10M0N(A1, B, NA2, Z);
  input A1, B, NA2;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(B_bar, B);
    and SMC_I2(OUT0, A1_bar, B_bar);
    and SMC_I3(OUT1, B_bar, NA2);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc NA2 --> Z
    (NA2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI21B10M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:06:55 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21B10M1N(A1, B, NA2, Z);
  input A1, B, NA2;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(B_bar, B);
    and SMC_I2(OUT0, A1_bar, B_bar);
    and SMC_I3(OUT1, B_bar, NA2);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc NA2 --> Z
    (NA2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI21B10M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:02:31 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21B10M2N(A1, B, NA2, Z);
  input A1, B, NA2;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(B_bar, B);
    and SMC_I2(OUT0, A1_bar, B_bar);
    and SMC_I3(OUT1, B_bar, NA2);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc NA2 --> Z
    (NA2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI21B10M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:09:36 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21B10M4N(A1, B, NA2, Z);
  input A1, B, NA2;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(B_bar, B);
    and SMC_I2(OUT0, A1_bar, B_bar);
    and SMC_I3(OUT1, B_bar, NA2);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc NA2 --> Z
    (NA2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI21B10M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:02:28 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21B20M0N(B, NA1, NA2, Z);
  input B, NA1, NA2;
  output Z;

    not SMC_I0(B_bar, B);
    and SMC_I1(OUT0, B_bar, NA2);
    and SMC_I2(OUT1, B_bar, NA1);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc NA1 --> Z
    (NA1 => Z) = (1.0, 1.0);

    // arc NA2 --> Z
    (NA2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI21B20M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:03:30 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21B20M1N(B, NA1, NA2, Z);
  input B, NA1, NA2;
  output Z;

    not SMC_I0(B_bar, B);
    and SMC_I1(OUT0, B_bar, NA2);
    and SMC_I2(OUT1, B_bar, NA1);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc NA1 --> Z
    (NA1 => Z) = (1.0, 1.0);

    // arc NA2 --> Z
    (NA2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI21B20M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:04:56 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21B20M2N(B, NA1, NA2, Z);
  input B, NA1, NA2;
  output Z;

    not SMC_I0(B_bar, B);
    and SMC_I1(OUT0, B_bar, NA2);
    and SMC_I2(OUT1, B_bar, NA1);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc NA1 --> Z
    (NA1 => Z) = (1.0, 1.0);

    // arc NA2 --> Z
    (NA2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI21B20M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:07:10 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21B20M4N(B, NA1, NA2, Z);
  input B, NA1, NA2;
  output Z;

    not SMC_I0(B_bar, B);
    and SMC_I1(OUT0, B_bar, NA2);
    and SMC_I2(OUT1, B_bar, NA1);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc NA1 --> Z
    (NA1 => Z) = (1.0, 1.0);

    // arc NA2 --> Z
    (NA2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI21B20M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:08:33 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21M0N(A1, A2, B, Z);
  input A1, A2, B;
  output Z;

    not SMC_I0(A2_bar, A2);
    not SMC_I1(B_bar, B);
    and SMC_I2(OUT0, A2_bar, B_bar);
    not SMC_I3(A1_bar, A1);
    and SMC_I4(OUT1, A1_bar, B_bar);
    or SMC_I5(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI21M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:04:14 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21M1N(A1, A2, B, Z);
  input A1, A2, B;
  output Z;

    not SMC_I0(A2_bar, A2);
    not SMC_I1(B_bar, B);
    and SMC_I2(OUT0, A2_bar, B_bar);
    not SMC_I3(A1_bar, A1);
    and SMC_I4(OUT1, A1_bar, B_bar);
    or SMC_I5(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI21M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:10:37 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21M2N(A1, A2, B, Z);
  input A1, A2, B;
  output Z;

    not SMC_I0(A2_bar, A2);
    not SMC_I1(B_bar, B);
    and SMC_I2(OUT0, A2_bar, B_bar);
    not SMC_I3(A1_bar, A1);
    and SMC_I4(OUT1, A1_bar, B_bar);
    or SMC_I5(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI21M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:02:47 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21M3N(A1, A2, B, Z);
  input A1, A2, B;
  output Z;

    not SMC_I0(A2_bar, A2);
    not SMC_I1(B_bar, B);
    and SMC_I2(OUT0, A2_bar, B_bar);
    not SMC_I3(A1_bar, A1);
    and SMC_I4(OUT1, A1_bar, B_bar);
    or SMC_I5(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI21M3N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:02:45 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21M4N(A1, A2, B, Z);
  input A1, A2, B;
  output Z;

    not SMC_I0(A2_bar, A2);
    not SMC_I1(B_bar, B);
    and SMC_I2(OUT0, A2_bar, B_bar);
    not SMC_I3(A1_bar, A1);
    and SMC_I4(OUT1, A1_bar, B_bar);
    or SMC_I5(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI21M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:05:12 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21M6N(A1, A2, B, Z);
  input A1, A2, B;
  output Z;

    not SMC_I0(A2_bar, A2);
    not SMC_I1(B_bar, B);
    and SMC_I2(OUT0, A2_bar, B_bar);
    not SMC_I3(A1_bar, A1);
    and SMC_I4(OUT1, A1_bar, B_bar);
    or SMC_I5(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI21M6N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:07:26 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21M8N(A1, A2, B, Z);
  input A1, A2, B;
  output Z;

    not SMC_I0(A2_bar, A2);
    not SMC_I1(B_bar, B);
    and SMC_I2(OUT0, A2_bar, B_bar);
    not SMC_I3(A1_bar, A1);
    and SMC_I4(OUT1, A1_bar, B_bar);
    or SMC_I5(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI21M8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:07:53 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI221M0N ( Z, A1, A2, B1, B2, C );
   input A1, A2, B1, B2, C;
   output Z;
      AOI221M0N_UDP5(Z, A1, A2, B1, B2, C);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI221M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:08:49 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI221M1N ( Z, A1, A2, B1, B2, C );
   input A1, A2, B1, B2, C;
   output Z;
      AOI221M0N_UDP5(Z, A1, A2, B1, B2, C);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI221M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:05:26 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI221M2N ( Z, A1, A2, B1, B2, C );
   input A1, A2, B1, B2, C;
   output Z;
      AOI221M0N_UDP5(Z, A1, A2, B1, B2, C);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI221M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:07:41 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI221M4N ( Z, A1, A2, B1, B2, C );
   input A1, A2, B1, B2, C;
   output Z;
      AOI221M0N_UDP5(Z, A1, A2, B1, B2, C);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI221M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:03:02 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI222M0N ( Z, A1, A2, B1, B2, C1, C2 );
   input A1, A2, B1, B2, C1, C2;
   output Z;
      AOI222M0N_UDP6(Z, A1, A2, B1, B2, C1, C2);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);

    // arc C1 --> Z
    (C1 => Z) = (1.0, 1.0);

    // arc C2 --> Z
    (C2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI222M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:02:59 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI222M1N ( Z, A1, A2, B1, B2, C1, C2 );
   input A1, A2, B1, B2, C1, C2;
   output Z;
      AOI222M0N_UDP6(Z, A1, A2, B1, B2, C1, C2);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);

    // arc C1 --> Z
    (C1 => Z) = (1.0, 1.0);

    // arc C2 --> Z
    (C2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI222M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:08:08 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI222M2N ( Z, A1, A2, B1, B2, C1, C2 );
   input A1, A2, B1, B2, C1, C2;
   output Z;
      AOI222M0N_UDP6(Z, A1, A2, B1, B2, C1, C2);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);

    // arc C1 --> Z
    (C1 => Z) = (1.0, 1.0);

    // arc C2 --> Z
    (C2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI222M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:09:03 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI222M4N ( Z, A1, A2, B1, B2, C1, C2 );
   input A1, A2, B1, B2, C1, C2;
   output Z;
      AOI222M0N_UDP6(Z, A1, A2, B1, B2, C1, C2);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);

    // arc C1 --> Z
    (C1 => Z) = (1.0, 1.0);

    // arc C2 --> Z
    (C2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI222M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:05:42 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI22B20M0N(B1, B2, NA1, NA2, Z);
  input B1, B2, NA1, NA2;
  output Z;

    not SMC_I0(B1_bar, B1);
    and SMC_I1(OUT0, B1_bar, NA1);
    not SMC_I2(B2_bar, B2);
    and SMC_I3(OUT1, B2_bar, NA1);
    and SMC_I4(OUT2, B1_bar, NA2);
    and SMC_I5(OUT3, B2_bar, NA2);
    or SMC_I6(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);

    // arc NA1 --> Z
    (NA1 => Z) = (1.0, 1.0);

    // arc NA2 --> Z
    (NA2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI22B20M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:07:56 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI22B20M1N(B1, B2, NA1, NA2, Z);
  input B1, B2, NA1, NA2;
  output Z;

    not SMC_I0(B1_bar, B1);
    and SMC_I1(OUT0, B1_bar, NA1);
    not SMC_I2(B2_bar, B2);
    and SMC_I3(OUT1, B2_bar, NA1);
    and SMC_I4(OUT2, B1_bar, NA2);
    and SMC_I5(OUT3, B2_bar, NA2);
    or SMC_I6(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);

    // arc NA1 --> Z
    (NA1 => Z) = (1.0, 1.0);

    // arc NA2 --> Z
    (NA2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI22B20M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:06:32 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI22B20M2N(B1, B2, NA1, NA2, Z);
  input B1, B2, NA1, NA2;
  output Z;

    not SMC_I0(B1_bar, B1);
    and SMC_I1(OUT0, B1_bar, NA1);
    not SMC_I2(B2_bar, B2);
    and SMC_I3(OUT1, B2_bar, NA1);
    and SMC_I4(OUT2, B1_bar, NA2);
    and SMC_I5(OUT3, B2_bar, NA2);
    or SMC_I6(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);

    // arc NA1 --> Z
    (NA1 => Z) = (1.0, 1.0);

    // arc NA2 --> Z
    (NA2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI22B20M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:09:05 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI22B20M4N(B1, B2, NA1, NA2, Z);
  input B1, B2, NA1, NA2;
  output Z;

    not SMC_I0(B1_bar, B1);
    and SMC_I1(OUT0, B1_bar, NA1);
    not SMC_I2(B2_bar, B2);
    and SMC_I3(OUT1, B2_bar, NA1);
    and SMC_I4(OUT2, B1_bar, NA2);
    and SMC_I5(OUT3, B2_bar, NA2);
    or SMC_I6(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);

    // arc NA1 --> Z
    (NA1 => Z) = (1.0, 1.0);

    // arc NA2 --> Z
    (NA2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI22B20M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:10:41 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI22M0N(A1, A2, B1, B2, Z);
  input A1, A2, B1, B2;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(B1_bar, B1);
    and SMC_I2(OUT0, A1_bar, B1_bar);
    not SMC_I3(A2_bar, A2);
    and SMC_I4(OUT1, A2_bar, B1_bar);
    not SMC_I5(B2_bar, B2);
    and SMC_I6(OUT2, A2_bar, B2_bar);
    and SMC_I7(OUT3, A1_bar, B2_bar);
    or SMC_I8(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI22M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:06:04 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI22M1N(A1, A2, B1, B2, Z);
  input A1, A2, B1, B2;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(B1_bar, B1);
    and SMC_I2(OUT0, A1_bar, B1_bar);
    not SMC_I3(A2_bar, A2);
    and SMC_I4(OUT1, A2_bar, B1_bar);
    not SMC_I5(B2_bar, B2);
    and SMC_I6(OUT2, A2_bar, B2_bar);
    and SMC_I7(OUT3, A1_bar, B2_bar);
    or SMC_I8(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI22M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:04:27 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI22M2N(A1, A2, B1, B2, Z);
  input A1, A2, B1, B2;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(B1_bar, B1);
    and SMC_I2(OUT0, A1_bar, B1_bar);
    not SMC_I3(A2_bar, A2);
    and SMC_I4(OUT1, A2_bar, B1_bar);
    not SMC_I5(B2_bar, B2);
    and SMC_I6(OUT2, A2_bar, B2_bar);
    and SMC_I7(OUT3, A1_bar, B2_bar);
    or SMC_I8(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI22M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:08:18 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI22M4N(A1, A2, B1, B2, Z);
  input A1, A2, B1, B2;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(B1_bar, B1);
    and SMC_I2(OUT0, A1_bar, B1_bar);
    not SMC_I3(A2_bar, A2);
    and SMC_I4(OUT1, A2_bar, B1_bar);
    not SMC_I5(B2_bar, B2);
    and SMC_I6(OUT2, A2_bar, B2_bar);
    and SMC_I7(OUT3, A1_bar, B2_bar);
    or SMC_I8(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI22M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:09:37 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI31M0N(A1, A2, A3, B, Z);
  input A1, A2, A3, B;
  output Z;

    not SMC_I0(A3_bar, A3);
    not SMC_I1(B_bar, B);
    and SMC_I2(OUT0, A3_bar, B_bar);
    not SMC_I3(A2_bar, A2);
    and SMC_I4(OUT1, A2_bar, B_bar);
    not SMC_I5(A1_bar, A1);
    and SMC_I6(OUT2, A1_bar, B_bar);
    or SMC_I7(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc A3 --> Z
    (A3 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI31M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:03:42 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI31M1N(A1, A2, A3, B, Z);
  input A1, A2, A3, B;
  output Z;

    not SMC_I0(A3_bar, A3);
    not SMC_I1(B_bar, B);
    and SMC_I2(OUT0, A3_bar, B_bar);
    not SMC_I3(A2_bar, A2);
    and SMC_I4(OUT1, A2_bar, B_bar);
    not SMC_I5(A1_bar, A1);
    and SMC_I6(OUT2, A1_bar, B_bar);
    or SMC_I7(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc A3 --> Z
    (A3 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI31M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:08:39 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI31M2N(A1, A2, A3, B, Z);
  input A1, A2, A3, B;
  output Z;

    not SMC_I0(A3_bar, A3);
    not SMC_I1(B_bar, B);
    and SMC_I2(OUT0, A3_bar, B_bar);
    not SMC_I3(A2_bar, A2);
    and SMC_I4(OUT1, A2_bar, B_bar);
    not SMC_I5(A1_bar, A1);
    and SMC_I6(OUT2, A1_bar, B_bar);
    or SMC_I7(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc A3 --> Z
    (A3 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI31M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:03:30 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI31M4N(A1, A2, A3, B, Z);
  input A1, A2, A3, B;
  output Z;

    not SMC_I0(A3_bar, A3);
    not SMC_I1(B_bar, B);
    and SMC_I2(OUT0, A3_bar, B_bar);
    not SMC_I3(A2_bar, A2);
    and SMC_I4(OUT1, A2_bar, B_bar);
    not SMC_I5(A1_bar, A1);
    and SMC_I6(OUT2, A1_bar, B_bar);
    or SMC_I7(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc A3 --> Z
    (A3 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI31M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:09:06 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI32M0N(A1, A2, A3, B1, B2, Z);
  input A1, A2, A3, B1, B2;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(B2_bar, B2);
    and SMC_I2(OUT0, A1_bar, B2_bar);
    not SMC_I3(A3_bar, A3);
    not SMC_I4(B1_bar, B1);
    and SMC_I5(OUT1, A3_bar, B1_bar);
    and SMC_I6(OUT2, A1_bar, B1_bar);
    and SMC_I7(OUT3, A3_bar, B2_bar);
    not SMC_I8(A2_bar, A2);
    and SMC_I9(OUT4, A2_bar, B1_bar);
    and SMC_I10(OUT5, A2_bar, B2_bar);
    or SMC_I11(Z, OUT0, OUT1, OUT2, OUT3, OUT4, OUT5);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc A3 --> Z
    (A3 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI32M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:06:34 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI32M1N(A1, A2, A3, B1, B2, Z);
  input A1, A2, A3, B1, B2;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(B2_bar, B2);
    and SMC_I2(OUT0, A1_bar, B2_bar);
    not SMC_I3(A3_bar, A3);
    not SMC_I4(B1_bar, B1);
    and SMC_I5(OUT1, A3_bar, B1_bar);
    and SMC_I6(OUT2, A1_bar, B1_bar);
    and SMC_I7(OUT3, A3_bar, B2_bar);
    not SMC_I8(A2_bar, A2);
    and SMC_I9(OUT4, A2_bar, B1_bar);
    and SMC_I10(OUT5, A2_bar, B2_bar);
    or SMC_I11(Z, OUT0, OUT1, OUT2, OUT3, OUT4, OUT5);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc A3 --> Z
    (A3 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI32M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:06:00 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI32M2N(A1, A2, A3, B1, B2, Z);
  input A1, A2, A3, B1, B2;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(B2_bar, B2);
    and SMC_I2(OUT0, A1_bar, B2_bar);
    not SMC_I3(A3_bar, A3);
    not SMC_I4(B1_bar, B1);
    and SMC_I5(OUT1, A3_bar, B1_bar);
    and SMC_I6(OUT2, A1_bar, B1_bar);
    and SMC_I7(OUT3, A3_bar, B2_bar);
    not SMC_I8(A2_bar, A2);
    and SMC_I9(OUT4, A2_bar, B1_bar);
    and SMC_I10(OUT5, A2_bar, B2_bar);
    or SMC_I11(Z, OUT0, OUT1, OUT2, OUT3, OUT4, OUT5);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc A3 --> Z
    (A3 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI32M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:03:35 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI32M4N(A1, A2, A3, B1, B2, Z);
  input A1, A2, A3, B1, B2;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(B2_bar, B2);
    and SMC_I2(OUT0, A1_bar, B2_bar);
    not SMC_I3(A3_bar, A3);
    not SMC_I4(B1_bar, B1);
    and SMC_I5(OUT1, A3_bar, B1_bar);
    and SMC_I6(OUT2, A1_bar, B1_bar);
    and SMC_I7(OUT3, A3_bar, B2_bar);
    not SMC_I8(A2_bar, A2);
    and SMC_I9(OUT4, A2_bar, B1_bar);
    and SMC_I10(OUT5, A2_bar, B2_bar);
    or SMC_I11(Z, OUT0, OUT1, OUT2, OUT3, OUT4, OUT5);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc A3 --> Z
    (A3 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI32M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:08:51 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI33M0N(A1, A2, A3, B1, B2, B3, Z);
  input A1, A2, A3, B1, B2, B3;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(B1_bar, B1);
    and SMC_I2(OUT0, A1_bar, B1_bar);
    not SMC_I3(A3_bar, A3);
    not SMC_I4(B3_bar, B3);
    and SMC_I5(OUT1, A3_bar, B3_bar);
    and SMC_I6(OUT2, A1_bar, B3_bar);
    not SMC_I7(A2_bar, A2);
    and SMC_I8(OUT3, A2_bar, B1_bar);
    not SMC_I9(B2_bar, B2);
    and SMC_I10(OUT4, A3_bar, B2_bar);
    and SMC_I11(OUT5, A2_bar, B2_bar);
    and SMC_I12(OUT6, A2_bar, B3_bar);
    and SMC_I13(OUT7, A3_bar, B1_bar);
    and SMC_I14(OUT8, A1_bar, B2_bar);
    or SMC_I15(OUTSUB0, OUT0, OUT1, OUT2, OUT3, OUT4, OUT5, OUT6, OUT7);
    or SMC_I16(OUTSUB1, OUT8);
    or SMC_I17(Z, OUTSUB0, OUTSUB1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc A3 --> Z
    (A3 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);

    // arc B3 --> Z
    (B3 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI33M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:09:48 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI33M1N(A1, A2, A3, B1, B2, B3, Z);
  input A1, A2, A3, B1, B2, B3;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(B1_bar, B1);
    and SMC_I2(OUT0, A1_bar, B1_bar);
    not SMC_I3(A3_bar, A3);
    not SMC_I4(B3_bar, B3);
    and SMC_I5(OUT1, A3_bar, B3_bar);
    and SMC_I6(OUT2, A1_bar, B3_bar);
    not SMC_I7(A2_bar, A2);
    and SMC_I8(OUT3, A2_bar, B1_bar);
    not SMC_I9(B2_bar, B2);
    and SMC_I10(OUT4, A3_bar, B2_bar);
    and SMC_I11(OUT5, A2_bar, B2_bar);
    and SMC_I12(OUT6, A2_bar, B3_bar);
    and SMC_I13(OUT7, A3_bar, B1_bar);
    and SMC_I14(OUT8, A1_bar, B2_bar);
    or SMC_I15(OUTSUB0, OUT0, OUT1, OUT2, OUT3, OUT4, OUT5, OUT6, OUT7);
    or SMC_I16(OUTSUB1, OUT8);
    or SMC_I17(Z, OUTSUB0, OUTSUB1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc A3 --> Z
    (A3 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);

    // arc B3 --> Z
    (B3 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI33M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:08:41 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI33M2N(A1, A2, A3, B1, B2, B3, Z);
  input A1, A2, A3, B1, B2, B3;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(B1_bar, B1);
    and SMC_I2(OUT0, A1_bar, B1_bar);
    not SMC_I3(A3_bar, A3);
    not SMC_I4(B3_bar, B3);
    and SMC_I5(OUT1, A3_bar, B3_bar);
    and SMC_I6(OUT2, A1_bar, B3_bar);
    not SMC_I7(A2_bar, A2);
    and SMC_I8(OUT3, A2_bar, B1_bar);
    not SMC_I9(B2_bar, B2);
    and SMC_I10(OUT4, A3_bar, B2_bar);
    and SMC_I11(OUT5, A2_bar, B2_bar);
    and SMC_I12(OUT6, A2_bar, B3_bar);
    and SMC_I13(OUT7, A3_bar, B1_bar);
    and SMC_I14(OUT8, A1_bar, B2_bar);
    or SMC_I15(OUTSUB0, OUT0, OUT1, OUT2, OUT3, OUT4, OUT5, OUT6, OUT7);
    or SMC_I16(OUTSUB1, OUT8);
    or SMC_I17(Z, OUTSUB0, OUTSUB1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc A3 --> Z
    (A3 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);

    // arc B3 --> Z
    (B3 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI33M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:09:35 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI33M4N(A1, A2, A3, B1, B2, B3, Z);
  input A1, A2, A3, B1, B2, B3;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(B1_bar, B1);
    and SMC_I2(OUT0, A1_bar, B1_bar);
    not SMC_I3(A3_bar, A3);
    not SMC_I4(B3_bar, B3);
    and SMC_I5(OUT1, A3_bar, B3_bar);
    and SMC_I6(OUT2, A1_bar, B3_bar);
    not SMC_I7(A2_bar, A2);
    and SMC_I8(OUT3, A2_bar, B1_bar);
    not SMC_I9(B2_bar, B2);
    and SMC_I10(OUT4, A3_bar, B2_bar);
    and SMC_I11(OUT5, A2_bar, B2_bar);
    and SMC_I12(OUT6, A2_bar, B3_bar);
    and SMC_I13(OUT7, A3_bar, B1_bar);
    and SMC_I14(OUT8, A1_bar, B2_bar);
    or SMC_I15(OUTSUB0, OUT0, OUT1, OUT2, OUT3, OUT4, OUT5, OUT6, OUT7);
    or SMC_I16(OUTSUB1, OUT8);
    or SMC_I17(Z, OUTSUB0, OUTSUB1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc A3 --> Z
    (A3 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);

    // arc B3 --> Z
    (B3 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // AOI33M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:07:18 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BEM1N(M0, M1, M2, OA1, OA2, Z);
  input M0, M1, M2;
  output OA1, OA2, Z;

    and SMC_I0(OUT0, M0, M1);
    not SMC_I1(M2_bar, M2);
    buf SMC_I2(OUT1, M2_bar);
    or SMC_I3(OA1, OUT0, OUT1);

    not SMC_I4(M0_bar, M0);
    not SMC_I5(M1_bar, M1);
    and SMC_I6(OUT2, M0_bar, M1_bar);
    buf SMC_I7(OUT3, M2);
    or SMC_I8(OA2, OUT2, OUT3);

    xnor SMC_I9(Z, M0, M1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc M0 --> OA1
    (M0 => OA1) = (1.0, 1.0);

    // arc M0 --> OA2
    (M0 => OA2) = (1.0, 1.0);

    // arc M0 --> Z
    if (M2===1'b0) 
        ( posedge M0 => ( Z +: M0 ) ) = (1.0, 1.0);
    if (M2===1'b0) 
        ( negedge M0 => ( Z +: M0 ) ) = (1.0, 1.0);
    if (M2===1'b1) 
        ( posedge M0 => ( Z +: M0 ) ) = (1.0, 1.0);
    if (M2===1'b1) 
        ( negedge M0 => ( Z +: M0 ) ) = (1.0, 1.0);
    ifnone
        ( posedge M0 => ( Z +: M0 ) ) = (1.0, 1.0);
        ( negedge M0 => ( Z +: M0 ) ) = (1.0, 1.0);

    // arc M1 --> OA1
    (M1 => OA1) = (1.0, 1.0);

    // arc M1 --> OA2
    (M1 => OA2) = (1.0, 1.0);

    // arc M1 --> Z
    if (M2===1'b0) 
        ( posedge M1 => ( Z +: M1 ) ) = (1.0, 1.0);
    if (M2===1'b0) 
        ( negedge M1 => ( Z +: M1 ) ) = (1.0, 1.0);
    if (M2===1'b1) 
        ( posedge M1 => ( Z +: M1 ) ) = (1.0, 1.0);
    if (M2===1'b1) 
        ( negedge M1 => ( Z +: M1 ) ) = (1.0, 1.0);
    ifnone
        ( posedge M1 => ( Z +: M1 ) ) = (1.0, 1.0);
        ( negedge M1 => ( Z +: M1 ) ) = (1.0, 1.0);

    // arc M2 --> OA1
    if (M0===1'b0 && M1===1'b0) 
        (M2 => OA1) = (1.0, 1.0);
    if (M0===1'b0 && M1===1'b1) 
        (M2 => OA1) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b0) 
        (M2 => OA1) = (1.0, 1.0);
    ifnone
        (M2 => OA1) = (1.0, 1.0);

    // arc M2 --> OA2
    if (M0===1'b0 && M1===1'b1) 
        (M2 => OA2) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b0) 
        (M2 => OA2) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b1) 
        (M2 => OA2) = (1.0, 1.0);
    ifnone
        (M2 => OA2) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // BEM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:06:47 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BEM2N(M0, M1, M2, OA1, OA2, Z);
  input M0, M1, M2;
  output OA1, OA2, Z;

    and SMC_I0(OUT0, M0, M1);
    not SMC_I1(M2_bar, M2);
    buf SMC_I2(OUT1, M2_bar);
    or SMC_I3(OA1, OUT0, OUT1);

    not SMC_I4(M0_bar, M0);
    not SMC_I5(M1_bar, M1);
    and SMC_I6(OUT2, M0_bar, M1_bar);
    buf SMC_I7(OUT3, M2);
    or SMC_I8(OA2, OUT2, OUT3);

    xnor SMC_I9(Z, M0, M1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc M0 --> OA1
    (M0 => OA1) = (1.0, 1.0);

    // arc M0 --> OA2
    (M0 => OA2) = (1.0, 1.0);

    // arc M0 --> Z
    if (M2===1'b0) 
        ( posedge M0 => ( Z +: M0 ) ) = (1.0, 1.0);
    if (M2===1'b0) 
        ( negedge M0 => ( Z +: M0 ) ) = (1.0, 1.0);
    if (M2===1'b1) 
        ( posedge M0 => ( Z +: M0 ) ) = (1.0, 1.0);
    if (M2===1'b1) 
        ( negedge M0 => ( Z +: M0 ) ) = (1.0, 1.0);
    ifnone
        ( posedge M0 => ( Z +: M0 ) ) = (1.0, 1.0);
        ( negedge M0 => ( Z +: M0 ) ) = (1.0, 1.0);

    // arc M1 --> OA1
    (M1 => OA1) = (1.0, 1.0);

    // arc M1 --> OA2
    (M1 => OA2) = (1.0, 1.0);

    // arc M1 --> Z
    if (M2===1'b0) 
        ( posedge M1 => ( Z +: M1 ) ) = (1.0, 1.0);
    if (M2===1'b0) 
        ( negedge M1 => ( Z +: M1 ) ) = (1.0, 1.0);
    if (M2===1'b1) 
        ( posedge M1 => ( Z +: M1 ) ) = (1.0, 1.0);
    if (M2===1'b1) 
        ( negedge M1 => ( Z +: M1 ) ) = (1.0, 1.0);
    ifnone
        ( posedge M1 => ( Z +: M1 ) ) = (1.0, 1.0);
        ( negedge M1 => ( Z +: M1 ) ) = (1.0, 1.0);

    // arc M2 --> OA1
    if (M0===1'b0 && M1===1'b0) 
        (M2 => OA1) = (1.0, 1.0);
    if (M0===1'b0 && M1===1'b1) 
        (M2 => OA1) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b0) 
        (M2 => OA1) = (1.0, 1.0);
    ifnone
        (M2 => OA1) = (1.0, 1.0);

    // arc M2 --> OA2
    if (M0===1'b0 && M1===1'b1) 
        (M2 => OA2) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b0) 
        (M2 => OA2) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b1) 
        (M2 => OA2) = (1.0, 1.0);
    ifnone
        (M2 => OA2) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // BEM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:05:03 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BEM4N(M0, M1, M2, OA1, OA2, Z);
  input M0, M1, M2;
  output OA1, OA2, Z;

    and SMC_I0(OUT0, M0, M1);
    not SMC_I1(M2_bar, M2);
    buf SMC_I2(OUT1, M2_bar);
    or SMC_I3(OA1, OUT0, OUT1);

    not SMC_I4(M0_bar, M0);
    not SMC_I5(M1_bar, M1);
    and SMC_I6(OUT2, M0_bar, M1_bar);
    buf SMC_I7(OUT3, M2);
    or SMC_I8(OA2, OUT2, OUT3);

    xnor SMC_I9(Z, M0, M1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc M0 --> OA1
    (M0 => OA1) = (1.0, 1.0);

    // arc M0 --> OA2
    (M0 => OA2) = (1.0, 1.0);

    // arc M0 --> Z
    if (M2===1'b0) 
        ( posedge M0 => ( Z +: M0 ) ) = (1.0, 1.0);
    if (M2===1'b0) 
        ( negedge M0 => ( Z +: M0 ) ) = (1.0, 1.0);
    if (M2===1'b1) 
        ( posedge M0 => ( Z +: M0 ) ) = (1.0, 1.0);
    if (M2===1'b1) 
        ( negedge M0 => ( Z +: M0 ) ) = (1.0, 1.0);
    ifnone
        ( posedge M0 => ( Z +: M0 ) ) = (1.0, 1.0);
        ( negedge M0 => ( Z +: M0 ) ) = (1.0, 1.0);

    // arc M1 --> OA1
    (M1 => OA1) = (1.0, 1.0);

    // arc M1 --> OA2
    (M1 => OA2) = (1.0, 1.0);

    // arc M1 --> Z
    if (M2===1'b0) 
        ( posedge M1 => ( Z +: M1 ) ) = (1.0, 1.0);
    if (M2===1'b0) 
        ( negedge M1 => ( Z +: M1 ) ) = (1.0, 1.0);
    if (M2===1'b1) 
        ( posedge M1 => ( Z +: M1 ) ) = (1.0, 1.0);
    if (M2===1'b1) 
        ( negedge M1 => ( Z +: M1 ) ) = (1.0, 1.0);
    ifnone
        ( posedge M1 => ( Z +: M1 ) ) = (1.0, 1.0);
        ( negedge M1 => ( Z +: M1 ) ) = (1.0, 1.0);

    // arc M2 --> OA1
    if (M0===1'b0 && M1===1'b0) 
        (M2 => OA1) = (1.0, 1.0);
    if (M0===1'b0 && M1===1'b1) 
        (M2 => OA1) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b0) 
        (M2 => OA1) = (1.0, 1.0);
    ifnone
        (M2 => OA1) = (1.0, 1.0);

    // arc M2 --> OA2
    if (M0===1'b0 && M1===1'b1) 
        (M2 => OA2) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b0) 
        (M2 => OA2) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b1) 
        (M2 => OA2) = (1.0, 1.0);
    ifnone
        (M2 => OA2) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // BEM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:11:28 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module BEMXBM2N ( PB, M0, M1, OA1, OA2, Z );
   input M0, M1, OA1, OA2, Z;
   output PB;
      BEMXBM2N_UDP5(PB, M0, M1, OA1, OA2, Z);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc M0 --> PB
    if (M1===1'b0) 
        ( posedge M0 => ( PB +: M0 ) ) = (1.0, 1.0);
    if (M1===1'b0) 
        ( negedge M0 => ( PB +: M0 ) ) = (1.0, 1.0);
    if (M1===1'b1) 
        ( posedge M0 => ( PB +: M0 ) ) = (1.0, 1.0);
    if (M1===1'b1) 
        ( negedge M0 => ( PB +: M0 ) ) = (1.0, 1.0);
    ifnone
        ( posedge M0 => ( PB +: M0 ) ) = (1.0, 1.0);
        ( negedge M0 => ( PB +: M0 ) ) = (1.0, 1.0);

    // arc M1 --> PB
    if (M0===1'b0) 
        ( posedge M1 => ( PB +: M1 ) ) = (1.0, 1.0);
    if (M0===1'b0) 
        ( negedge M1 => ( PB +: M1 ) ) = (1.0, 1.0);
    if (M0===1'b1) 
        ( posedge M1 => ( PB +: M1 ) ) = (1.0, 1.0);
    if (M0===1'b1) 
        ( negedge M1 => ( PB +: M1 ) ) = (1.0, 1.0);
    ifnone
        ( posedge M1 => ( PB +: M1 ) ) = (1.0, 1.0);
        ( negedge M1 => ( PB +: M1 ) ) = (1.0, 1.0);

    // arc OA1 --> PB
    if (M0===1'b0 && M1===1'b1 && OA2===1'b0 && Z===1'b0) 
        (OA1 => PB) = (1.0, 1.0);
    if (M0===1'b0 && M1===1'b1 && OA2===1'b1 && Z===1'b0) 
        (OA1 => PB) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b0 && OA2===1'b0 && Z===1'b1) 
        (OA1 => PB) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b0 && OA2===1'b1 && Z===1'b1) 
        (OA1 => PB) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b1 && OA2===1'b0 && Z===1'b0) 
        (OA1 => PB) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b1 && OA2===1'b0 && Z===1'b1) 
        (OA1 => PB) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b1 && OA2===1'b1 && Z===1'b0) 
        (OA1 => PB) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b1 && OA2===1'b1 && Z===1'b1) 
        (OA1 => PB) = (1.0, 1.0);
    ifnone
        (OA1 => PB) = (1.0, 1.0);

    // arc OA2 --> PB
    if (M0===1'b0 && M1===1'b0 && OA1===1'b0 && Z===1'b0) 
        (OA2 => PB) = (1.0, 1.0);
    if (M0===1'b0 && M1===1'b0 && OA1===1'b0 && Z===1'b1) 
        (OA2 => PB) = (1.0, 1.0);
    if (M0===1'b0 && M1===1'b0 && OA1===1'b1 && Z===1'b0) 
        (OA2 => PB) = (1.0, 1.0);
    if (M0===1'b0 && M1===1'b0 && OA1===1'b1 && Z===1'b1) 
        (OA2 => PB) = (1.0, 1.0);
    if (M0===1'b0 && M1===1'b1 && OA1===1'b0 && Z===1'b1) 
        (OA2 => PB) = (1.0, 1.0);
    if (M0===1'b0 && M1===1'b1 && OA1===1'b1 && Z===1'b1) 
        (OA2 => PB) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b0 && OA1===1'b0 && Z===1'b0) 
        (OA2 => PB) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b0 && OA1===1'b1 && Z===1'b0) 
        (OA2 => PB) = (1.0, 1.0);
    ifnone
        (OA2 => PB) = (1.0, 1.0);

    // arc Z --> PB
    if (M0===1'b0 && M1===1'b1 && OA1===1'b0 && OA2===1'b1) 
        (Z => PB) = (1.0, 1.0);
    if (M0===1'b0 && M1===1'b1 && OA1===1'b1 && OA2===1'b0) 
        (Z => PB) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b0 && OA1===1'b0 && OA2===1'b1) 
        (Z => PB) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b0 && OA1===1'b1 && OA2===1'b0) 
        (Z => PB) = (1.0, 1.0);
    ifnone
        ( posedge Z => ( PB +: Z ) ) = (1.0, 1.0);
        ( negedge Z => ( PB +: Z ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // BEMXBM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:09:32 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module BEMXBM4N ( PB, M0, M1, OA1, OA2, Z );
   input M0, M1, OA1, OA2, Z;
   output PB;
      BEMXBM2N_UDP5(PB, M0, M1, OA1, OA2, Z);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc M0 --> PB
    if (M1===1'b0) 
        ( posedge M0 => ( PB +: M0 ) ) = (1.0, 1.0);
    if (M1===1'b0) 
        ( negedge M0 => ( PB +: M0 ) ) = (1.0, 1.0);
    if (M1===1'b1) 
        ( posedge M0 => ( PB +: M0 ) ) = (1.0, 1.0);
    if (M1===1'b1) 
        ( negedge M0 => ( PB +: M0 ) ) = (1.0, 1.0);
    ifnone
        ( posedge M0 => ( PB +: M0 ) ) = (1.0, 1.0);
        ( negedge M0 => ( PB +: M0 ) ) = (1.0, 1.0);

    // arc M1 --> PB
    if (M0===1'b0) 
        ( posedge M1 => ( PB +: M1 ) ) = (1.0, 1.0);
    if (M0===1'b0) 
        ( negedge M1 => ( PB +: M1 ) ) = (1.0, 1.0);
    if (M0===1'b1) 
        ( posedge M1 => ( PB +: M1 ) ) = (1.0, 1.0);
    if (M0===1'b1) 
        ( negedge M1 => ( PB +: M1 ) ) = (1.0, 1.0);
    ifnone
        ( posedge M1 => ( PB +: M1 ) ) = (1.0, 1.0);
        ( negedge M1 => ( PB +: M1 ) ) = (1.0, 1.0);

    // arc OA1 --> PB
    if (M0===1'b0 && M1===1'b1 && OA2===1'b0 && Z===1'b0) 
        (OA1 => PB) = (1.0, 1.0);
    if (M0===1'b0 && M1===1'b1 && OA2===1'b1 && Z===1'b0) 
        (OA1 => PB) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b0 && OA2===1'b0 && Z===1'b1) 
        (OA1 => PB) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b0 && OA2===1'b1 && Z===1'b1) 
        (OA1 => PB) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b1 && OA2===1'b0 && Z===1'b0) 
        (OA1 => PB) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b1 && OA2===1'b0 && Z===1'b1) 
        (OA1 => PB) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b1 && OA2===1'b1 && Z===1'b0) 
        (OA1 => PB) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b1 && OA2===1'b1 && Z===1'b1) 
        (OA1 => PB) = (1.0, 1.0);
    ifnone
        (OA1 => PB) = (1.0, 1.0);

    // arc OA2 --> PB
    if (M0===1'b0 && M1===1'b0 && OA1===1'b0 && Z===1'b0) 
        (OA2 => PB) = (1.0, 1.0);
    if (M0===1'b0 && M1===1'b0 && OA1===1'b0 && Z===1'b1) 
        (OA2 => PB) = (1.0, 1.0);
    if (M0===1'b0 && M1===1'b0 && OA1===1'b1 && Z===1'b0) 
        (OA2 => PB) = (1.0, 1.0);
    if (M0===1'b0 && M1===1'b0 && OA1===1'b1 && Z===1'b1) 
        (OA2 => PB) = (1.0, 1.0);
    if (M0===1'b0 && M1===1'b1 && OA1===1'b0 && Z===1'b1) 
        (OA2 => PB) = (1.0, 1.0);
    if (M0===1'b0 && M1===1'b1 && OA1===1'b1 && Z===1'b1) 
        (OA2 => PB) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b0 && OA1===1'b0 && Z===1'b0) 
        (OA2 => PB) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b0 && OA1===1'b1 && Z===1'b0) 
        (OA2 => PB) = (1.0, 1.0);
    ifnone
        (OA2 => PB) = (1.0, 1.0);

    // arc Z --> PB
    if (M0===1'b0 && M1===1'b1 && OA1===1'b0 && OA2===1'b1) 
        (Z => PB) = (1.0, 1.0);
    if (M0===1'b0 && M1===1'b1 && OA1===1'b1 && OA2===1'b0) 
        (Z => PB) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b0 && OA1===1'b0 && OA2===1'b1) 
        (Z => PB) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b0 && OA1===1'b1 && OA2===1'b0) 
        (Z => PB) = (1.0, 1.0);
    ifnone
        ( posedge Z => ( PB +: Z ) ) = (1.0, 1.0);
        ( negedge Z => ( PB +: Z ) ) = (1.0, 1.0);


   endspecify

  `endif // functional //
endmodule     // BEMXBM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:10:38 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module BEMXM2N ( P, M0, M1, OA1, OA2, Z );
   input M0, M1, OA1, OA2, Z;
   output P;
      BEMXM2N_UDP5(P, M0, M1, OA1, OA2, Z);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc M0 --> P
    if (M1===1'b0) 
        ( posedge M0 => ( P +: M0 ) ) = (1.0, 1.0);
    if (M1===1'b0) 
        ( negedge M0 => ( P +: M0 ) ) = (1.0, 1.0);
    if (M1===1'b1) 
        ( posedge M0 => ( P +: M0 ) ) = (1.0, 1.0);
    if (M1===1'b1) 
        ( negedge M0 => ( P +: M0 ) ) = (1.0, 1.0);
    ifnone
        ( posedge M0 => ( P +: M0 ) ) = (1.0, 1.0);
        ( negedge M0 => ( P +: M0 ) ) = (1.0, 1.0);

    // arc M1 --> P
    if (M0===1'b0) 
        ( posedge M1 => ( P +: M1 ) ) = (1.0, 1.0);
    if (M0===1'b0) 
        ( negedge M1 => ( P +: M1 ) ) = (1.0, 1.0);
    if (M0===1'b1) 
        ( posedge M1 => ( P +: M1 ) ) = (1.0, 1.0);
    if (M0===1'b1) 
        ( negedge M1 => ( P +: M1 ) ) = (1.0, 1.0);
    ifnone
        ( posedge M1 => ( P +: M1 ) ) = (1.0, 1.0);
        ( negedge M1 => ( P +: M1 ) ) = (1.0, 1.0);

    // arc OA1 --> P
    if (M0===1'b0 && M1===1'b1 && OA2===1'b0 && Z===1'b0) 
        (OA1 => P) = (1.0, 1.0);
    if (M0===1'b0 && M1===1'b1 && OA2===1'b1 && Z===1'b0) 
        (OA1 => P) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b0 && OA2===1'b0 && Z===1'b1) 
        (OA1 => P) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b0 && OA2===1'b1 && Z===1'b1) 
        (OA1 => P) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b1 && OA2===1'b0 && Z===1'b0) 
        (OA1 => P) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b1 && OA2===1'b0 && Z===1'b1) 
        (OA1 => P) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b1 && OA2===1'b1 && Z===1'b0) 
        (OA1 => P) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b1 && OA2===1'b1 && Z===1'b1) 
        (OA1 => P) = (1.0, 1.0);
    ifnone
        (OA1 => P) = (1.0, 1.0);

    // arc OA2 --> P
    if (M0===1'b0 && M1===1'b0 && OA1===1'b0 && Z===1'b0) 
        (OA2 => P) = (1.0, 1.0);
    if (M0===1'b0 && M1===1'b0 && OA1===1'b0 && Z===1'b1) 
        (OA2 => P) = (1.0, 1.0);
    if (M0===1'b0 && M1===1'b0 && OA1===1'b1 && Z===1'b0) 
        (OA2 => P) = (1.0, 1.0);
    if (M0===1'b0 && M1===1'b0 && OA1===1'b1 && Z===1'b1) 
        (OA2 => P) = (1.0, 1.0);
    if (M0===1'b0 && M1===1'b1 && OA1===1'b0 && Z===1'b1) 
        (OA2 => P) = (1.0, 1.0);
    if (M0===1'b0 && M1===1'b1 && OA1===1'b1 && Z===1'b1) 
        (OA2 => P) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b0 && OA1===1'b0 && Z===1'b0) 
        (OA2 => P) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b0 && OA1===1'b1 && Z===1'b0) 
        (OA2 => P) = (1.0, 1.0);
    ifnone
        (OA2 => P) = (1.0, 1.0);

    // arc Z --> P
    if (M0===1'b0 && M1===1'b1 && OA1===1'b0 && OA2===1'b1) 
        (Z => P) = (1.0, 1.0);
    if (M0===1'b0 && M1===1'b1 && OA1===1'b1 && OA2===1'b0) 
        (Z => P) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b0 && OA1===1'b0 && OA2===1'b1) 
        (Z => P) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b0 && OA1===1'b1 && OA2===1'b0) 
        (Z => P) = (1.0, 1.0);
    ifnone
        ( posedge Z => ( P +: Z ) ) = (1.0, 1.0);
        ( negedge Z => ( P +: Z ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // BEMXM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:04:41 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module BEMXM4N ( P, M0, M1, OA1, OA2, Z );
   input M0, M1, OA1, OA2, Z;
   output P;
      BEMXM2N_UDP5(P, M0, M1, OA1, OA2, Z);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc M0 --> P
    if (M1===1'b0) 
        ( posedge M0 => ( P +: M0 ) ) = (1.0, 1.0);
    if (M1===1'b0) 
        ( negedge M0 => ( P +: M0 ) ) = (1.0, 1.0);
    if (M1===1'b1) 
        ( posedge M0 => ( P +: M0 ) ) = (1.0, 1.0);
    if (M1===1'b1) 
        ( negedge M0 => ( P +: M0 ) ) = (1.0, 1.0);
    ifnone
        ( posedge M0 => ( P +: M0 ) ) = (1.0, 1.0);
        ( negedge M0 => ( P +: M0 ) ) = (1.0, 1.0);

    // arc M1 --> P
    if (M0===1'b0) 
        ( posedge M1 => ( P +: M1 ) ) = (1.0, 1.0);
    if (M0===1'b0) 
        ( negedge M1 => ( P +: M1 ) ) = (1.0, 1.0);
    if (M0===1'b1) 
        ( posedge M1 => ( P +: M1 ) ) = (1.0, 1.0);
    if (M0===1'b1) 
        ( negedge M1 => ( P +: M1 ) ) = (1.0, 1.0);
    ifnone
        ( posedge M1 => ( P +: M1 ) ) = (1.0, 1.0);
        ( negedge M1 => ( P +: M1 ) ) = (1.0, 1.0);

    // arc OA1 --> P
    if (M0===1'b0 && M1===1'b1 && OA2===1'b0 && Z===1'b0) 
        (OA1 => P) = (1.0, 1.0);
    if (M0===1'b0 && M1===1'b1 && OA2===1'b1 && Z===1'b0) 
        (OA1 => P) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b0 && OA2===1'b0 && Z===1'b1) 
        (OA1 => P) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b0 && OA2===1'b1 && Z===1'b1) 
        (OA1 => P) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b1 && OA2===1'b0 && Z===1'b0) 
        (OA1 => P) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b1 && OA2===1'b0 && Z===1'b1) 
        (OA1 => P) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b1 && OA2===1'b1 && Z===1'b0) 
        (OA1 => P) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b1 && OA2===1'b1 && Z===1'b1) 
        (OA1 => P) = (1.0, 1.0);
    ifnone
        (OA1 => P) = (1.0, 1.0);

    // arc OA2 --> P
    if (M0===1'b0 && M1===1'b0 && OA1===1'b0 && Z===1'b0) 
        (OA2 => P) = (1.0, 1.0);
    if (M0===1'b0 && M1===1'b0 && OA1===1'b0 && Z===1'b1) 
        (OA2 => P) = (1.0, 1.0);
    if (M0===1'b0 && M1===1'b0 && OA1===1'b1 && Z===1'b0) 
        (OA2 => P) = (1.0, 1.0);
    if (M0===1'b0 && M1===1'b0 && OA1===1'b1 && Z===1'b1) 
        (OA2 => P) = (1.0, 1.0);
    if (M0===1'b0 && M1===1'b1 && OA1===1'b0 && Z===1'b1) 
        (OA2 => P) = (1.0, 1.0);
    if (M0===1'b0 && M1===1'b1 && OA1===1'b1 && Z===1'b1) 
        (OA2 => P) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b0 && OA1===1'b0 && Z===1'b0) 
        (OA2 => P) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b0 && OA1===1'b1 && Z===1'b0) 
        (OA2 => P) = (1.0, 1.0);
    ifnone
        (OA2 => P) = (1.0, 1.0);

    // arc Z --> P
    if (M0===1'b0 && M1===1'b1 && OA1===1'b0 && OA2===1'b1) 
        (Z => P) = (1.0, 1.0);
    if (M0===1'b0 && M1===1'b1 && OA1===1'b1 && OA2===1'b0) 
        (Z => P) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b0 && OA1===1'b0 && OA2===1'b1) 
        (Z => P) = (1.0, 1.0);
    if (M0===1'b1 && M1===1'b0 && OA1===1'b1 && OA2===1'b0) 
        (Z => P) = (1.0, 1.0);
    ifnone
        ( posedge Z => ( P +: Z ) ) = (1.0, 1.0);
        ( negedge Z => ( P +: Z ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // BEMXM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:04:39 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BHDM1N(Z);
  inout Z;

  // Busholder.
  wire io_wire;

  buf(weak0,weak1) SMC_I0(Z, io_wire);
  buf              SMC_I1(io_wire, Z);

  `ifdef functional // functional //

  `else // functional //

  specify




  endspecify

  `endif // functional //
endmodule     // BHDM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:04:38 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFM10N(A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // BUFM10N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:06:48 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFM12N(A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // BUFM12N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:09:21 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFM14N(A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // BUFM14N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:06:14 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFM16N(A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // BUFM16N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:08:28 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFM18N(A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // BUFM18N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:10:54 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFM20N(A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // BUFM20N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:03:49 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFM2N(A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // BUFM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:06:49 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFM3N(A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // BUFM3N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:06:14 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFM4N(A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // BUFM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:09:22 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFM5N(A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // BUFM5N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:05:34 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFM6N(A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // BUFM6N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:08:29 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFM8N(A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // BUFM8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:10:55 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFTM0N(A, E, Z);
  input A, E;
  output Z;

    buf SMC_I0(SMC_DIN0, A);

    not SMC_I1(SMC_ZEN0, E);


    bufif0 SMC_I2(Z, SMC_DIN0, SMC_ZEN0);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc E --> Z
    (E => Z) = (1.0,
        1.0,
        1.0,
        1.0,
        1.0,
        1.0);



  endspecify

  `endif // functional //
endmodule     // BUFTM0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:08:56 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFTM12N(A, E, Z);
  input A, E;
  output Z;

    buf SMC_I0(SMC_DIN0, A);

    not SMC_I1(SMC_ZEN0, E);


    bufif0 SMC_I2(Z, SMC_DIN0, SMC_ZEN0);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc E --> Z
    (E => Z) = (1.0,
        1.0,
        1.0,
        1.0,
        1.0,
        1.0);



  endspecify

  `endif // functional //
endmodule     // BUFTM12N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:09:52 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFTM16N(A, E, Z);
  input A, E;
  output Z;

    buf SMC_I0(SMC_DIN0, A);

    not SMC_I1(SMC_ZEN0, E);


    bufif0 SMC_I2(Z, SMC_DIN0, SMC_ZEN0);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc E --> Z
    (E => Z) = (1.0,
        1.0,
        1.0,
        1.0,
        1.0,
        1.0);



  endspecify

  `endif // functional //
endmodule     // BUFTM16N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:03:48 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFTM1N(A, E, Z);
  input A, E;
  output Z;

    buf SMC_I0(SMC_DIN0, A);

    not SMC_I1(SMC_ZEN0, E);


    bufif0 SMC_I2(Z, SMC_DIN0, SMC_ZEN0);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc E --> Z
    (E => Z) = (1.0,
        1.0,
        1.0,
        1.0,
        1.0,
        1.0);



  endspecify

  `endif // functional //
endmodule     // BUFTM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:03:50 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFTM20N(A, E, Z);
  input A, E;
  output Z;

    buf SMC_I0(SMC_DIN0, A);

    not SMC_I1(SMC_ZEN0, E);


    bufif0 SMC_I2(Z, SMC_DIN0, SMC_ZEN0);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc E --> Z
    (E => Z) = (1.0,
        1.0,
        1.0,
        1.0,
        1.0,
        1.0);



  endspecify

  `endif // functional //
endmodule     // BUFTM20N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:09:38 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFTM2N(A, E, Z);
  input A, E;
  output Z;

    buf SMC_I0(SMC_DIN0, A);

    not SMC_I1(SMC_ZEN0, E);


    bufif0 SMC_I2(Z, SMC_DIN0, SMC_ZEN0);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc E --> Z
    (E => Z) = (1.0,
        1.0,
        1.0,
        1.0,
        1.0,
        1.0);



  endspecify

  `endif // functional //
endmodule     // BUFTM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:08:45 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFTM3N(A, E, Z);
  input A, E;
  output Z;

    buf SMC_I0(SMC_DIN0, A);

    not SMC_I1(SMC_ZEN0, E);


    bufif0 SMC_I2(Z, SMC_DIN0, SMC_ZEN0);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc E --> Z
    (E => Z) = (1.0,
        1.0,
        1.0,
        1.0,
        1.0,
        1.0);



  endspecify

  `endif // functional //
endmodule     // BUFTM3N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:07:06 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFTM4N(A, E, Z);
  input A, E;
  output Z;

    buf SMC_I0(SMC_DIN0, A);

    not SMC_I1(SMC_ZEN0, E);


    bufif0 SMC_I2(Z, SMC_DIN0, SMC_ZEN0);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc E --> Z
    (E => Z) = (1.0,
        1.0,
        1.0,
        1.0,
        1.0,
        1.0);



  endspecify

  `endif // functional //
endmodule     // BUFTM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:06:31 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFTM6N(A, E, Z);
  input A, E;
  output Z;

    buf SMC_I0(SMC_DIN0, A);

    not SMC_I1(SMC_ZEN0, E);


    bufif0 SMC_I2(Z, SMC_DIN0, SMC_ZEN0);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc E --> Z
    (E => Z) = (1.0,
        1.0,
        1.0,
        1.0,
        1.0,
        1.0);



  endspecify

  `endif // functional //
endmodule     // BUFTM6N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:11:12 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFTM8N(A, E, Z);
  input A, E;
  output Z;

    buf SMC_I0(SMC_DIN0, A);

    not SMC_I1(SMC_ZEN0, E);


    bufif0 SMC_I2(Z, SMC_DIN0, SMC_ZEN0);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc E --> Z
    (E => Z) = (1.0,
        1.0,
        1.0,
        1.0,
        1.0,
        1.0);



  endspecify

  `endif // functional //
endmodule     // BUFTM8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:04:07 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKAN2M12N(A, B, Z);
  input A, B;
  output Z;

    and SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // CKAN2M12N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:08:47 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKAN2M2N(A, B, Z);
  input A, B;
  output Z;

    and SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // CKAN2M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:07:06 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKAN2M3N(A, B, Z);
  input A, B;
  output Z;

    and SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // CKAN2M3N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:09:40 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKAN2M4N(A, B, Z);
  input A, B;
  output Z;

    and SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // CKAN2M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:04:54 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKAN2M6N(A, B, Z);
  input A, B;
  output Z;

    and SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // CKAN2M6N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:06:33 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKAN2M8N(A, B, Z);
  input A, B;
  output Z;

    and SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // CKAN2M8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:11:15 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKBUFM12N(A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // CKBUFM12N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:09:15 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKBUFM16N(A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // CKBUFM16N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:10:12 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKBUFM1N(A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // CKBUFM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:04:08 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKBUFM20N(A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // CKBUFM20N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:04:11 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKBUFM24N(A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // CKBUFM24N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:04:11 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKBUFM2N(A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // CKBUFM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:07:11 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKBUFM32N(A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // CKBUFM32N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:09:44 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKBUFM3N(A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // CKBUFM3N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:04:56 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKBUFM40N(A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // CKBUFM40N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:08:50 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKBUFM4N(A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // CKBUFM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:07:15 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKBUFM6N(A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // CKBUFM6N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:11:17 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKBUFM8N(A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // CKBUFM8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:09:18 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKINVM12N(A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // CKINVM12N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:04:12 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKINVM16N(A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // CKINVM16N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:10:14 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKINVM1N(A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // CKINVM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:07:37 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKINVM20N(A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // CKINVM20N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:09:16 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKINVM24N(A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // CKINVM24N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:10:10 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKINVM2N(A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // CKINVM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:07:38 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKINVM32N(A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // CKINVM32N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:05:22 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKINVM3N(A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // CKINVM3N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:07:03 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKINVM40N(A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // CKINVM40N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:10:41 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKINVM4N(A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // CKINVM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:11:44 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKINVM6N(A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // CKINVM6N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:04:39 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKINVM8N(A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // CKINVM8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:09:18 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKMUX2M12N(A, B, S, Z);
  input A, B, S;
  output Z;

    not SMC_I0(S_bar, S);
    and SMC_I1(OUT0, A, S_bar);
    and SMC_I2(OUT1, B, S);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        (A => Z) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        (B => Z) = (1.0, 1.0);

    // arc S --> Z
     if ( S===1'b1 )
    ( posedge S => ( Z +: S ) ) = (1.0, 1.0);
     if ( S===1'b0 )
    ( negedge S => ( Z +: S ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // CKMUX2M12N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:09:45 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKMUX2M2N(A, B, S, Z);
  input A, B, S;
  output Z;

    not SMC_I0(S_bar, S);
    and SMC_I1(OUT0, A, S_bar);
    and SMC_I2(OUT1, B, S);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        (A => Z) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        (B => Z) = (1.0, 1.0);

    // arc S --> Z
     if ( S===1'b1 )
    ( posedge S => ( Z +: S ) ) = (1.0, 1.0);
     if ( S===1'b0 )
    ( negedge S => ( Z +: S ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // CKMUX2M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:10:11 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKMUX2M3N(A, B, S, Z);
  input A, B, S;
  output Z;

    not SMC_I0(S_bar, S);
    and SMC_I1(OUT0, A, S_bar);
    and SMC_I2(OUT1, B, S);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        (A => Z) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        (B => Z) = (1.0, 1.0);

    // arc S --> Z
     if ( S===1'b1 )
    ( posedge S => ( Z +: S ) ) = (1.0, 1.0);
     if ( S===1'b0 )
    ( negedge S => ( Z +: S ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // CKMUX2M3N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:05:24 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKMUX2M4N(A, B, S, Z);
  input A, B, S;
  output Z;

    not SMC_I0(S_bar, S);
    and SMC_I1(OUT0, A, S_bar);
    and SMC_I2(OUT1, B, S);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        (A => Z) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        (B => Z) = (1.0, 1.0);

    // arc S --> Z
     if ( S===1'b1 )
    ( posedge S => ( Z +: S ) ) = (1.0, 1.0);
     if ( S===1'b0 )
    ( negedge S => ( Z +: S ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // CKMUX2M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:07:51 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKMUX2M6N(A, B, S, Z);
  input A, B, S;
  output Z;

    not SMC_I0(S_bar, S);
    and SMC_I1(OUT0, A, S_bar);
    and SMC_I2(OUT1, B, S);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        (A => Z) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        (B => Z) = (1.0, 1.0);

    // arc S --> Z
     if ( S===1'b1 )
    ( posedge S => ( Z +: S ) ) = (1.0, 1.0);
     if ( S===1'b0 )
    ( negedge S => ( Z +: S ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // CKMUX2M6N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:04:38 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKMUX2M8N(A, B, S, Z);
  input A, B, S;
  output Z;

    not SMC_I0(S_bar, S);
    and SMC_I1(OUT0, A, S_bar);
    and SMC_I2(OUT1, B, S);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        (A => Z) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        (B => Z) = (1.0, 1.0);

    // arc S --> Z
     if ( S===1'b1 )
    ( posedge S => ( Z +: S ) ) = (1.0, 1.0);
     if ( S===1'b0 )
    ( negedge S => ( Z +: S ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // CKMUX2M8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:07:15 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKND2M12N(A, B, Z);
  input A, B;
  output Z;

    nand SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // CKND2M12N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:11:59 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKND2M2N(A, B, Z);
  input A, B;
  output Z;

    nand SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // CKND2M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:10:13 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKND2M4N(A, B, Z);
  input A, B;
  output Z;

    nand SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // CKND2M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:10:01 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKND2M8N(A, B, Z);
  input A, B;
  output Z;

    nand SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // CKND2M8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:09:35 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKXOR2M12N(A, B, Z);
  input A, B;
  output Z;

    xor SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
     if ( A===1'b1 )
    ( posedge A => ( Z +: A ) ) = (1.0, 1.0);
     if ( A===1'b0 )
    ( negedge A => ( Z +: A ) ) = (1.0, 1.0);

    // arc B --> Z
     if ( B===1'b1 )
    ( posedge B => ( Z +: B ) ) = (1.0, 1.0);
     if ( B===1'b0 )
    ( negedge B => ( Z +: B ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // CKXOR2M12N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:04:41 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKXOR2M1N(A, B, Z);
  input A, B;
  output Z;

    xor SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (  A => Z ) = (1.0, 1.0);
     if ( A===1'b1 )
    ( posedge A => ( Z +: A ) ) = (1.0, 1.0);
     if ( A===1'b0 )
    ( negedge A => ( Z +: A ) ) = (1.0, 1.0);

    // arc B --> Z
     if ( B===1'b1 )
    ( posedge B => ( Z +: B ) ) = (1.0, 1.0);
     if ( B===1'b0 )
    ( negedge B => ( Z +: B ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // CKXOR2M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:10:43 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKXOR2M2N(A, B, Z);
  input A, B;
  output Z;

    xor SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
     if ( A===1'b1 )
    ( posedge A => ( Z +: A ) ) = (1.0, 1.0);
     if ( A===1'b0 )
    ( negedge A => ( Z +: A ) ) = (1.0, 1.0);

    // arc B --> Z
     if ( B===1'b1 )
    ( posedge B => ( Z +: B ) ) = (1.0, 1.0);
     if ( B===1'b0 )
    ( negedge B => ( Z +: B ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // CKXOR2M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:04:58 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKXOR2M4N(A, B, Z);
  input A, B;
  output Z;

    xor SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
     if ( A===1'b1 )
    ( posedge A => ( Z +: A ) ) = (1.0, 1.0);
     if ( A===1'b0 )
    ( negedge A => ( Z +: A ) ) = (1.0, 1.0);

    // arc B --> Z
     if ( B===1'b1 )
    ( posedge B => ( Z +: B ) ) = (1.0, 1.0);
     if ( B===1'b0 )
    ( negedge B => ( Z +: B ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // CKXOR2M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:05:41 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKXOR2M8N(A, B, Z);
  input A, B;
  output Z;

    xor SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
     if ( A===1'b1 )
    ( posedge A => ( Z +: A ) ) = (1.0, 1.0);
     if ( A===1'b0 )
    ( negedge A => ( Z +: A ) ) = (1.0, 1.0);

    // arc B --> Z
     if ( B===1'b1 )
    ( posedge B => ( Z +: B ) ) = (1.0, 1.0);
     if ( B===1'b0 )
    ( negedge B => ( Z +: B ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // CKXOR2M8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:07:42 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DEL1M1N(A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // DEL1M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:07:07 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DEL1M4N(A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // DEL1M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:12:05 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DEL2M1N(A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // DEL2M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:05:00 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DEL2M4N(A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // DEL2M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:09:48 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DEL3M1N(A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // DEL3M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:09:21 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DEL3M4N(A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // DEL3M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:10:15 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DEL4M1N(A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // DEL4M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:10:23 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DEL4M4N(A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // DEL4M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:04:49 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFEM0N(D, E, CK, Q, QB);
  input D, E, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, D, SMC_IQ, E);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I6(shcheckCKDlh, E);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: E )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: E )) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // setup D-hl CK-lh (E)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (E)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // hold D-hl CK-lh (E)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (E)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFEM0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:07:34 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFEM1N(D, E, CK, Q, QB);
  input D, E, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, D, SMC_IQ, E);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I6(shcheckCKDlh, E);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: E )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: E )) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // setup D-hl CK-lh (E)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (E)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // hold D-hl CK-lh (E)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (E)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFEM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:08:07 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFEM2N(D, E, CK, Q, QB);
  input D, E, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, D, SMC_IQ, E);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I6(shcheckCKDlh, E);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: E )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: E )) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // setup D-hl CK-lh (E)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (E)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // hold D-hl CK-lh (E)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (E)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFEM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:05:52 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFEM4N(D, E, CK, Q, QB);
  input D, E, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, D, SMC_IQ, E);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I6(shcheckCKDlh, E);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: E )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: E )) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // setup D-hl CK-lh (E)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (E)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // hold D-hl CK-lh (E)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (E)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFEM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:10:42 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFEQBM0N(D, E, CK, QB);
  input D, E, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, D, SMC_IQ, E);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(shcheckCKDlh, E);


  specify


    // arc CK --> QB
    (posedge CK => ( QB +: E )) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // setup D-hl CK-lh (E)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (E)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // hold D-hl CK-lh (E)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (E)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFEQBM0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:12:14 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFEQBM1N(D, E, CK, QB);
  input D, E, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, D, SMC_IQ, E);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(shcheckCKDlh, E);


  specify


    // arc CK --> QB
    (posedge CK => ( QB +: E )) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // setup D-hl CK-lh (E)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (E)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // hold D-hl CK-lh (E)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (E)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFEQBM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:09:48 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFEQBM2N(D, E, CK, QB);
  input D, E, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, D, SMC_IQ, E);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(shcheckCKDlh, E);


  specify


    // arc CK --> QB
    (posedge CK => ( QB +: E )) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // setup D-hl CK-lh (E)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (E)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // hold D-hl CK-lh (E)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (E)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFEQBM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:10:16 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFEQBM4N(D, E, CK, QB);
  input D, E, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, D, SMC_IQ, E);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(shcheckCKDlh, E);


  specify


    // arc CK --> QB
    (posedge CK => ( QB +: E )) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // setup D-hl CK-lh (E)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (E)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // hold D-hl CK-lh (E)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (E)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFEQBM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:11:12 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFEZRM0N(D, E, RB, CK, Q, QB);
  input D, E, RB, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    DFEZRM0N_UDP__OUT__ SMC_I1(SMC_NS_IN, D, E, SMC_IQ, RB);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I6(shcheckCKDlh, E, RB);

    buf SMC_I7(shcheckCKElh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup E-hl CK-lh (RB)
    $setup(negedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // setup E-lh CK-lh (RB)
    $setup(posedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (E&RB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (E&RB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup RB-hl CK-lh ()
    $setup(negedge RB, posedge CK, 1.0, notifier);

    // setup RB-lh CK-lh ()
    $setup(posedge RB, posedge CK, 1.0, notifier);

    // hold E-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        negedge E &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // hold E-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        posedge E &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (E&RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (E&RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold RB-hl CK-lh ()
    $hold(posedge CK, negedge RB, 1.0, notifier);

    // hold RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFEZRM0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:05:08 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFEZRM1N(D, E, RB, CK, Q, QB);
  input D, E, RB, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    DFEZRM0N_UDP__OUT__ SMC_I1(SMC_NS_IN, D, E, SMC_IQ, RB);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I6(shcheckCKDlh, E, RB);

    buf SMC_I7(shcheckCKElh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup E-hl CK-lh (RB)
    $setup(negedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // setup E-lh CK-lh (RB)
    $setup(posedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (E&RB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (E&RB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup RB-hl CK-lh ()
    $setup(negedge RB, posedge CK, 1.0, notifier);

    // setup RB-lh CK-lh ()
    $setup(posedge RB, posedge CK, 1.0, notifier);

    // hold E-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        negedge E &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // hold E-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        posedge E &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (E&RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (E&RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold RB-hl CK-lh ()
    $hold(posedge CK, negedge RB, 1.0, notifier);

    // hold RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFEZRM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:05:11 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFEZRM2N(D, E, RB, CK, Q, QB);
  input D, E, RB, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    DFEZRM0N_UDP__OUT__ SMC_I1(SMC_NS_IN, D, E, SMC_IQ, RB);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I6(shcheckCKDlh, E, RB);

    buf SMC_I7(shcheckCKElh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup E-hl CK-lh (RB)
    $setup(negedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // setup E-lh CK-lh (RB)
    $setup(posedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (E&RB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (E&RB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup RB-hl CK-lh ()
    $setup(negedge RB, posedge CK, 1.0, notifier);

    // setup RB-lh CK-lh ()
    $setup(posedge RB, posedge CK, 1.0, notifier);

    // hold E-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        negedge E &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // hold E-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        posedge E &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (E&RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (E&RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold RB-hl CK-lh ()
    $hold(posedge CK, negedge RB, 1.0, notifier);

    // hold RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFEZRM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:05:11 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFEZRM4N(D, E, RB, CK, Q, QB);
  input D, E, RB, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    DFEZRM0N_UDP__OUT__ SMC_I1(SMC_NS_IN, D, E, SMC_IQ, RB);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I6(shcheckCKDlh, E, RB);

    buf SMC_I7(shcheckCKElh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup E-hl CK-lh (RB)
    $setup(negedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // setup E-lh CK-lh (RB)
    $setup(posedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (E&RB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (E&RB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup RB-hl CK-lh ()
    $setup(negedge RB, posedge CK, 1.0, notifier);

    // setup RB-lh CK-lh ()
    $setup(posedge RB, posedge CK, 1.0, notifier);

    // hold E-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        negedge E &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // hold E-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        posedge E &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (E&RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (E&RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold RB-hl CK-lh ()
    $hold(posedge CK, negedge RB, 1.0, notifier);

    // hold RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFEZRM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:05:11 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFM0N(D, CK, Q, QB);
  input D, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh ()
    $setup(posedge D, posedge CK, 1.0, notifier);

    // setup D-hl CK-lh ()
    $setup(negedge D, posedge CK, 1.0, notifier);

    // hold D-lh CK-lh ()
    $hold(posedge CK, posedge D, 1.0, notifier);

    // hold D-hl CK-lh ()
    $hold(posedge CK, negedge D, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFM0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:08:12 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFM1N(D, CK, Q, QB);
  input D, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh ()
    $setup(posedge D, posedge CK, 1.0, notifier);

    // setup D-hl CK-lh ()
    $setup(negedge D, posedge CK, 1.0, notifier);

    // hold D-lh CK-lh ()
    $hold(posedge CK, posedge D, 1.0, notifier);

    // hold D-hl CK-lh ()
    $hold(posedge CK, negedge D, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:09:55 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFM2N(D, CK, Q, QB);
  input D, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh ()
    $setup(posedge D, posedge CK, 1.0, notifier);

    // setup D-hl CK-lh ()
    $setup(negedge D, posedge CK, 1.0, notifier);

    // hold D-lh CK-lh ()
    $hold(posedge CK, posedge D, 1.0, notifier);

    // hold D-hl CK-lh ()
    $hold(posedge CK, negedge D, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:05:56 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFM4N(D, CK, Q, QB);
  input D, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh ()
    $setup(posedge D, posedge CK, 1.0, notifier);

    // setup D-hl CK-lh ()
    $setup(negedge D, posedge CK, 1.0, notifier);

    // hold D-lh CK-lh ()
    $hold(posedge CK, posedge D, 1.0, notifier);

    // hold D-hl CK-lh ()
    $hold(posedge CK, negedge D, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:07:41 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQBM0N(D, CK, QB);
  input D, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh ()
    $setup(negedge D, posedge CK, 1.0, notifier);

    // setup D-lh CK-lh ()
    $setup(posedge D, posedge CK, 1.0, notifier);

    // hold D-hl CK-lh ()
    $hold(posedge CK, negedge D, 1.0, notifier);

    // hold D-lh CK-lh ()
    $hold(posedge CK, posedge D, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQBM0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:12:18 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQBM1N(D, CK, QB);
  input D, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh ()
    $setup(negedge D, posedge CK, 1.0, notifier);

    // setup D-lh CK-lh ()
    $setup(posedge D, posedge CK, 1.0, notifier);

    // hold D-hl CK-lh ()
    $hold(posedge CK, negedge D, 1.0, notifier);

    // hold D-lh CK-lh ()
    $hold(posedge CK, posedge D, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQBM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:10:47 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQBM2N(D, CK, QB);
  input D, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh ()
    $setup(negedge D, posedge CK, 1.0, notifier);

    // setup D-lh CK-lh ()
    $setup(posedge D, posedge CK, 1.0, notifier);

    // hold D-hl CK-lh ()
    $hold(posedge CK, negedge D, 1.0, notifier);

    // hold D-lh CK-lh ()
    $hold(posedge CK, posedge D, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQBM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:10:23 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQBM4N(D, CK, QB);
  input D, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh ()
    $setup(negedge D, posedge CK, 1.0, notifier);

    // setup D-lh CK-lh ()
    $setup(posedge D, posedge CK, 1.0, notifier);

    // hold D-hl CK-lh ()
    $hold(posedge CK, negedge D, 1.0, notifier);

    // hold D-lh CK-lh ()
    $hold(posedge CK, posedge D, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQBM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:11:20 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQBRM0N(D, RB, CK, QB);
  input D, RB, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I4(shcheckCKDlh, RB);


  specify


    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (RB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (RB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 1.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQBRM0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:08:17 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQBRM1N(D, RB, CK, QB);
  input D, RB, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I4(shcheckCKDlh, RB);


  specify


    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (RB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (RB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 1.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQBRM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:06:05 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQBRM2N(D, RB, CK, QB);
  input D, RB, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I4(shcheckCKDlh, RB);


  specify


    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (RB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (RB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 1.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQBRM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:07:45 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQBRM4N(D, RB, CK, QB);
  input D, RB, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I4(shcheckCKDlh, RB);


  specify


    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (RB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (RB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 1.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQBRM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:10:48 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQM0N(D, CK, Q);
  input D, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh ()
    $setup(negedge D, posedge CK, 1.0, notifier);

    // setup D-lh CK-lh ()
    $setup(posedge D, posedge CK, 1.0, notifier);

    // hold D-hl CK-lh ()
    $hold(posedge CK, negedge D, 1.0, notifier);

    // hold D-lh CK-lh ()
    $hold(posedge CK, posedge D, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQM0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:09:55 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQM1N(D, CK, Q);
  input D, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh ()
    $setup(negedge D, posedge CK, 1.0, notifier);

    // setup D-lh CK-lh ()
    $setup(posedge D, posedge CK, 1.0, notifier);

    // hold D-hl CK-lh ()
    $hold(posedge CK, negedge D, 1.0, notifier);

    // hold D-lh CK-lh ()
    $hold(posedge CK, posedge D, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:12:21 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQM2N(D, CK, Q);
  input D, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh ()
    $setup(negedge D, posedge CK, 1.0, notifier);

    // setup D-lh CK-lh ()
    $setup(posedge D, posedge CK, 1.0, notifier);

    // hold D-hl CK-lh ()
    $hold(posedge CK, negedge D, 1.0, notifier);

    // hold D-lh CK-lh ()
    $hold(posedge CK, posedge D, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:11:17 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQM4N(D, CK, Q);
  input D, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh ()
    $setup(negedge D, posedge CK, 1.0, notifier);

    // setup D-lh CK-lh ()
    $setup(posedge D, posedge CK, 1.0, notifier);

    // hold D-hl CK-lh ()
    $hold(posedge CK, negedge D, 1.0, notifier);

    // hold D-lh CK-lh ()
    $hold(posedge CK, posedge D, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:10:22 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQRM0N(D, RB, CK, Q);
  input D, RB, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckCKDlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (RB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (RB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 1.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQRM0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:05:22 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQRM1N(D, RB, CK, Q);
  input D, RB, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckCKDlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (RB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (RB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 1.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQRM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:05:13 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQRM2N(D, RB, CK, Q);
  input D, RB, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckCKDlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (RB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (RB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 1.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQRM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:10:53 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQRM4N(D, RB, CK, Q);
  input D, RB, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckCKDlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (RB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (RB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 1.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQRM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:12:27 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQSM0N(D, SB, CK, Q);
  input D, SB, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //
    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(SB));

  `else // functional //
    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckCKDlh, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (SB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (SB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 1.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQSM0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:10:00 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQSM1N(D, SB, CK, Q);
  input D, SB, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //
    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(SB));

  `else // functional //
    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckCKDlh, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (SB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (SB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 1.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQSM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:10:28 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQSM2N(D, SB, CK, Q);
  input D, SB, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //
    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(SB));

  `else // functional //
    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckCKDlh, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (SB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (SB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 1.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQSM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:05:19 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQSM4N(D, SB, CK, Q);
  input D, SB, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //
    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(SB));

  `else // functional //
    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckCKDlh, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (SB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (SB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 1.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQSM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:05:24 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFRM0N(D, RB, CK, Q, QB);
  input D, RB, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(shcheckCKDlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (RB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (RB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 1.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFRM0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:05:25 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFRM1N(D, RB, CK, Q, QB);
  input D, RB, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(shcheckCKDlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (RB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (RB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 1.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFRM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:08:22 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFRM2N(D, RB, CK, Q, QB);
  input D, RB, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(shcheckCKDlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (RB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (RB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 1.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFRM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:07:48 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFRM4N(D, RB, CK, Q, QB);
  input D, RB, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(shcheckCKDlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (RB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (RB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 1.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFRM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:06:12 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFRSM0N(D, RB, SB, CK, Q, QB);
  input D, RB, SB, CK;
  output Q, QB;
  reg notifier;

    inv_clr0 SMC_I0(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ));

  `ifdef functional // functional //
    dff_p1 SMC_I2(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(SB));

  `else // functional //
    dff_p1 SMC_I2(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I6(shcheckCKDlh, RB, SB);

    buf SMC_I7(shcheckCKRBlh, SB);

    buf SMC_I8(shcheckCKSBlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (RB&SB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (RB&SB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SB-lh RB-lh ()
    $setup(posedge SB, posedge RB, 1.0, notifier);

    // hold D-hl CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SB-lh RB-lh ()
    $hold(posedge RB, posedge SB, 1.0, notifier);

    // recovery RB-lh CK-lh (SB)
    $recovery(posedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh (RB)
    $recovery(posedge SB &&& (shcheckCKSBlh === 1'b1),
        posedge CK &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // removal RB-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        posedge RB &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // removal SB-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSBlh === 1'b1),
        posedge SB &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFRSM0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:11:00 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFRSM1N(D, RB, SB, CK, Q, QB);
  input D, RB, SB, CK;
  output Q, QB;
  reg notifier;

    inv_clr0 SMC_I0(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ));

  `ifdef functional // functional //
    dff_p1 SMC_I2(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(SB));

  `else // functional //
    dff_p1 SMC_I2(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I6(shcheckCKDlh, RB, SB);

    buf SMC_I7(shcheckCKRBlh, SB);

    buf SMC_I8(shcheckCKSBlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (RB&SB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (RB&SB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SB-lh RB-lh ()
    $setup(posedge SB, posedge RB, 1.0, notifier);

    // hold D-hl CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SB-lh RB-lh ()
    $hold(posedge RB, posedge SB, 1.0, notifier);

    // recovery RB-lh CK-lh (SB)
    $recovery(posedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh (RB)
    $recovery(posedge SB &&& (shcheckCKSBlh === 1'b1),
        posedge CK &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // removal RB-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        posedge RB &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // removal SB-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSBlh === 1'b1),
        posedge SB &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFRSM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:12:28 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFRSM2N(D, RB, SB, CK, Q, QB);
  input D, RB, SB, CK;
  output Q, QB;
  reg notifier;

    inv_clr0 SMC_I0(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ));

  `ifdef functional // functional //
    dff_p1 SMC_I2(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(SB));

  `else // functional //
    dff_p1 SMC_I2(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I6(shcheckCKDlh, RB, SB);

    buf SMC_I7(shcheckCKRBlh, SB);

    buf SMC_I8(shcheckCKSBlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (RB&SB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (RB&SB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SB-lh RB-lh ()
    $setup(posedge SB, posedge RB, 1.0, notifier);

    // hold D-hl CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SB-lh RB-lh ()
    $hold(posedge RB, posedge SB, 1.0, notifier);

    // recovery RB-lh CK-lh (SB)
    $recovery(posedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh (RB)
    $recovery(posedge SB &&& (shcheckCKSBlh === 1'b1),
        posedge CK &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // removal RB-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        posedge RB &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // removal SB-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSBlh === 1'b1),
        posedge SB &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFRSM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:10:02 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFRSM4N(D, RB, SB, CK, Q, QB);
  input D, RB, SB, CK;
  output Q, QB;
  reg notifier;

    inv_clr0 SMC_I0(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ));

  `ifdef functional // functional //
    dff_p1 SMC_I2(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(SB));

  `else // functional //
    dff_p1 SMC_I2(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I6(shcheckCKDlh, RB, SB);

    buf SMC_I7(shcheckCKRBlh, SB);

    buf SMC_I8(shcheckCKSBlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (RB&SB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (RB&SB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SB-lh RB-lh ()
    $setup(posedge SB, posedge RB, 1.0, notifier);

    // hold D-hl CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SB-lh RB-lh ()
    $hold(posedge RB, posedge SB, 1.0, notifier);

    // recovery RB-lh CK-lh (SB)
    $recovery(posedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh (RB)
    $recovery(posedge SB &&& (shcheckCKSBlh === 1'b1),
        posedge CK &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // removal RB-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        posedge RB &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // removal SB-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSBlh === 1'b1),
        posedge SB &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFRSM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:10:30 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFSM0N(D, SB, CK, Q, QB);
  input D, SB, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(SB));

  `else // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(shcheckCKDlh, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (SB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (SB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 1.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFSM0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:11:26 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFSM1N(D, SB, CK, Q, QB);
  input D, SB, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(SB));

  `else // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(shcheckCKDlh, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (SB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (SB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 1.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFSM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:08:39 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFSM2N(D, SB, CK, Q, QB);
  input D, SB, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(SB));

  `else // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(shcheckCKDlh, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (SB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (SB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 1.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFSM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:06:23 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFSM4N(D, SB, CK, Q, QB);
  input D, SB, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(SB));

  `else // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(shcheckCKDlh, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (SB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (SB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 1.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFSM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:11:12 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFZRM0N(D, RB, CK, Q, QB);
  input D, RB, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    and SMC_I1(SMC_NS_IN, D, RB);


  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh ()
    $setup(negedge D, posedge CK, 1.0, notifier);

    // setup D-lh CK-lh ()
    $setup(posedge D, posedge CK, 1.0, notifier);

    // setup RB-hl CK-lh ()
    $setup(negedge RB, posedge CK, 1.0, notifier);

    // setup RB-lh CK-lh ()
    $setup(posedge RB, posedge CK, 1.0, notifier);

    // hold D-hl CK-lh ()
    $hold(posedge CK, negedge D, 1.0, notifier);

    // hold D-lh CK-lh ()
    $hold(posedge CK, posedge D, 1.0, notifier);

    // hold RB-hl CK-lh ()
    $hold(posedge CK, negedge RB, 1.0, notifier);

    // hold RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFZRM0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:08:05 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFZRM1N(D, RB, CK, Q, QB);
  input D, RB, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    and SMC_I1(SMC_NS_IN, D, RB);


  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh ()
    $setup(negedge D, posedge CK, 1.0, notifier);

    // setup D-lh CK-lh ()
    $setup(posedge D, posedge CK, 1.0, notifier);

    // setup RB-hl CK-lh ()
    $setup(negedge RB, posedge CK, 1.0, notifier);

    // setup RB-lh CK-lh ()
    $setup(posedge RB, posedge CK, 1.0, notifier);

    // hold D-hl CK-lh ()
    $hold(posedge CK, negedge D, 1.0, notifier);

    // hold D-lh CK-lh ()
    $hold(posedge CK, posedge D, 1.0, notifier);

    // hold RB-hl CK-lh ()
    $hold(posedge CK, negedge RB, 1.0, notifier);

    // hold RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFZRM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:12:46 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFZRM2N(D, RB, CK, Q, QB);
  input D, RB, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    and SMC_I1(SMC_NS_IN, D, RB);


  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh ()
    $setup(negedge D, posedge CK, 1.0, notifier);

    // setup D-lh CK-lh ()
    $setup(posedge D, posedge CK, 1.0, notifier);

    // setup RB-hl CK-lh ()
    $setup(negedge RB, posedge CK, 1.0, notifier);

    // setup RB-lh CK-lh ()
    $setup(posedge RB, posedge CK, 1.0, notifier);

    // hold D-hl CK-lh ()
    $hold(posedge CK, negedge D, 1.0, notifier);

    // hold D-lh CK-lh ()
    $hold(posedge CK, posedge D, 1.0, notifier);

    // hold RB-hl CK-lh ()
    $hold(posedge CK, negedge RB, 1.0, notifier);

    // hold RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFZRM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:10:19 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFZRM4N(D, RB, CK, Q, QB);
  input D, RB, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    and SMC_I1(SMC_NS_IN, D, RB);


  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh ()
    $setup(negedge D, posedge CK, 1.0, notifier);

    // setup D-lh CK-lh ()
    $setup(posedge D, posedge CK, 1.0, notifier);

    // setup RB-hl CK-lh ()
    $setup(negedge RB, posedge CK, 1.0, notifier);

    // setup RB-lh CK-lh ()
    $setup(posedge RB, posedge CK, 1.0, notifier);

    // hold D-hl CK-lh ()
    $hold(posedge CK, negedge D, 1.0, notifier);

    // hold D-lh CK-lh ()
    $hold(posedge CK, posedge D, 1.0, notifier);

    // hold RB-hl CK-lh ()
    $hold(posedge CK, negedge RB, 1.0, notifier);

    // hold RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFZRM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:11:42 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module HADFM0N ( CO, S, A, B, CI );
   input A, B, CI;
   output CO, S;
      ADFM0N_UDP3(CO, A, B, CI);
      ADFM0N_UDP4(S, A, B, CI);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO
    if (B===1'b0 && CI===1'b1) 
        (A => CO) = (1.0, 1.0);
    if (B===1'b1 && CI===1'b0) 
        (A => CO) = (1.0, 1.0);
    ifnone
        (A => CO) = (1.0, 1.0);

    // arc A --> S
    if (B===1'b0 && CI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && CI===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CI===1'b1) 
        (A => S) = (1.0, 1.0);
    ifnone
        ( posedge A => ( S +: A ) ) = (1.0, 1.0);
        ( negedge A => ( S +: A ) ) = (1.0, 1.0);

    // arc B --> CO
    if (A===1'b0 && CI===1'b1) 
        (B => CO) = (1.0, 1.0);
    if (A===1'b1 && CI===1'b0) 
        (B => CO) = (1.0, 1.0);
    ifnone
        (B => CO) = (1.0, 1.0);

    // arc B --> S
    if (A===1'b0 && CI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && CI===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CI===1'b1) 
        (B => S) = (1.0, 1.0);
    ifnone
        ( posedge B => ( S +: B ) ) = (1.0, 1.0);
        ( negedge B => ( S +: B ) ) = (1.0, 1.0);

    // arc CI --> CO
    if (A===1'b0 && B===1'b1) 
        (CI => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0) 
        (CI => CO) = (1.0, 1.0);
    ifnone
        (CI => CO) = (1.0, 1.0);

    // arc CI --> S
    if (A===1'b0 && B===1'b0) 
        (CI => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1) 
        (CI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0) 
        (CI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1) 
        (CI => S) = (1.0, 1.0);
    ifnone
        ( posedge CI => ( S +: CI ) ) = (1.0, 1.0);
        ( negedge CI => ( S +: CI ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // HADFM0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:05:43 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module HADFM1N ( CO, S, A, B, CI );
   input A, B, CI;
   output CO, S;
      ADFM0N_UDP3(CO, A, B, CI);
      ADFM0N_UDP4(S, A, B, CI);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO
    if (B===1'b0 && CI===1'b1) 
        (A => CO) = (1.0, 1.0);
    if (B===1'b1 && CI===1'b0) 
        (A => CO) = (1.0, 1.0);
    ifnone
        (A => CO) = (1.0, 1.0);

    // arc A --> S
    if (B===1'b0 && CI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && CI===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CI===1'b1) 
        (A => S) = (1.0, 1.0);
    ifnone
        ( posedge A => ( S +: A ) ) = (1.0, 1.0);
        ( negedge A => ( S +: A ) ) = (1.0, 1.0);

    // arc B --> CO
    if (A===1'b0 && CI===1'b1) 
        (B => CO) = (1.0, 1.0);
    if (A===1'b1 && CI===1'b0) 
        (B => CO) = (1.0, 1.0);
    ifnone
        (B => CO) = (1.0, 1.0);

    // arc B --> S
    if (A===1'b0 && CI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && CI===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CI===1'b1) 
        (B => S) = (1.0, 1.0);
    ifnone
        ( posedge B => ( S +: B ) ) = (1.0, 1.0);
        ( negedge B => ( S +: B ) ) = (1.0, 1.0);

    // arc CI --> CO
    if (A===1'b0 && B===1'b1) 
        (CI => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0) 
        (CI => CO) = (1.0, 1.0);
    ifnone
        (CI => CO) = (1.0, 1.0);

    // arc CI --> S
    if (A===1'b0 && B===1'b0) 
        (CI => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1) 
        (CI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0) 
        (CI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1) 
        (CI => S) = (1.0, 1.0);
    ifnone
        ( posedge CI => ( S +: CI ) ) = (1.0, 1.0);
        ( negedge CI => ( S +: CI ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // HADFM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:10:47 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module HADFM2N ( CO, S, A, B, CI );
   input A, B, CI;
   output CO, S;
      ADFM0N_UDP3(CO, A, B, CI);
      ADFM0N_UDP4(S, A, B, CI);
   
  `ifdef functional // functional //

  `else // functional //

 specify


    // arc A --> CO
    if (B===1'b0 && CI===1'b1) 
        (A => CO) = (1.0, 1.0);
    if (B===1'b1 && CI===1'b0) 
        (A => CO) = (1.0, 1.0);
    ifnone
        (A => CO) = (1.0, 1.0);

    // arc A --> S
    if (B===1'b0 && CI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && CI===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CI===1'b1) 
        (A => S) = (1.0, 1.0);
    ifnone
        ( posedge A => ( S +: A ) ) = (1.0, 1.0);
        ( negedge A => ( S +: A ) ) = (1.0, 1.0);

    // arc B --> CO
    if (A===1'b0 && CI===1'b1) 
        (B => CO) = (1.0, 1.0);
    if (A===1'b1 && CI===1'b0) 
        (B => CO) = (1.0, 1.0);
    ifnone
        (B => CO) = (1.0, 1.0);

    // arc B --> S
    if (A===1'b0 && CI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && CI===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CI===1'b1) 
        (B => S) = (1.0, 1.0);
    ifnone
        ( posedge B => ( S +: B ) ) = (1.0, 1.0);
        ( negedge B => ( S +: B ) ) = (1.0, 1.0);

    // arc CI --> CO
    if (A===1'b0 && B===1'b1) 
        (CI => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0) 
        (CI => CO) = (1.0, 1.0);
    ifnone
        (CI => CO) = (1.0, 1.0);

    // arc CI --> S
    if (A===1'b0 && B===1'b0) 
        (CI => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1) 
        (CI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0) 
        (CI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1) 
        (CI => S) = (1.0, 1.0);
    ifnone
        ( posedge CI => ( S +: CI ) ) = (1.0, 1.0);
        ( negedge CI => ( S +: CI ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // HADFM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:08:42 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module HADFM4N ( CO, S, A, B, CI );
   input A, B, CI;
   output CO, S;
      ADFM0N_UDP3(CO, A, B, CI);
      ADFM0N_UDP4(S, A, B, CI);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO
    if (B===1'b0 && CI===1'b1) 
        (A => CO) = (1.0, 1.0);
    if (B===1'b1 && CI===1'b0) 
        (A => CO) = (1.0, 1.0);
    ifnone
        (A => CO) = (1.0, 1.0);

    // arc A --> S
    if (B===1'b0 && CI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b0 && CI===1'b1) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CI===1'b0) 
        (A => S) = (1.0, 1.0);
    if (B===1'b1 && CI===1'b1) 
        (A => S) = (1.0, 1.0);
    ifnone
        ( posedge A => ( S +: A ) ) = (1.0, 1.0);
        ( negedge A => ( S +: A ) ) = (1.0, 1.0);

    // arc B --> CO
    if (A===1'b0 && CI===1'b1) 
        (B => CO) = (1.0, 1.0);
    if (A===1'b1 && CI===1'b0) 
        (B => CO) = (1.0, 1.0);
    ifnone
        (B => CO) = (1.0, 1.0);

    // arc B --> S
    if (A===1'b0 && CI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b0 && CI===1'b1) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CI===1'b0) 
        (B => S) = (1.0, 1.0);
    if (A===1'b1 && CI===1'b1) 
        (B => S) = (1.0, 1.0);
    ifnone
        ( posedge B => ( S +: B ) ) = (1.0, 1.0);
        ( negedge B => ( S +: B ) ) = (1.0, 1.0);

    // arc CI --> CO
    if (A===1'b0 && B===1'b1) 
        (CI => CO) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0) 
        (CI => CO) = (1.0, 1.0);
    ifnone
        (CI => CO) = (1.0, 1.0);

    // arc CI --> S
    if (A===1'b0 && B===1'b0) 
        (CI => S) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1) 
        (CI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0) 
        (CI => S) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1) 
        (CI => S) = (1.0, 1.0);
    ifnone
        ( posedge CI => ( S +: CI ) ) = (1.0, 1.0);
        ( negedge CI => ( S +: CI ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // HADFM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:08:10 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HDFCM1N(D, CKB, Q, QB);
  input D, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (1.0, 1.0);

    // arc CKB --> QB
    (negedge CKB => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CKB-hl ()
    $setup(posedge D, negedge CKB, 1.0, notifier);

    // setup D-hl CKB-hl ()
    $setup(negedge D, negedge CKB, 1.0, notifier);

    // hold D-lh CKB-hl ()
    $hold(negedge CKB, posedge D, 1.0, notifier);

    // hold D-hl CKB-hl ()
    $hold(negedge CKB, negedge D, 1.0, notifier);

    // mpw CKB-lh NS-lh ()
    $width(posedge CKB, 1.0, 0, notifier);

    // mpw CKB-hl NS-hl ()
    $width(negedge CKB, 1.0, 0, notifier);

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HDFCM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:05:39 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HDFCM2N(D, CKB, Q, QB);
  input D, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (1.0, 1.0);

    // arc CKB --> QB
    (negedge CKB => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CKB-hl ()
    $setup(posedge D, negedge CKB, 1.0, notifier);

    // setup D-hl CKB-hl ()
    $setup(negedge D, negedge CKB, 1.0, notifier);

    // hold D-lh CKB-hl ()
    $hold(negedge CKB, posedge D, 1.0, notifier);

    // hold D-hl CKB-hl ()
    $hold(negedge CKB, negedge D, 1.0, notifier);

    // mpw CKB-lh NS-lh ()
    $width(posedge CKB, 1.0, 0, notifier);

    // mpw CKB-hl NS-hl ()
    $width(negedge CKB, 1.0, 0, notifier);

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HDFCM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:05:41 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HDFCM4N(D, CKB, Q, QB);
  input D, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (1.0, 1.0);

    // arc CKB --> QB
    (negedge CKB => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CKB-hl ()
    $setup(posedge D, negedge CKB, 1.0, notifier);

    // setup D-hl CKB-hl ()
    $setup(negedge D, negedge CKB, 1.0, notifier);

    // hold D-lh CKB-hl ()
    $hold(negedge CKB, posedge D, 1.0, notifier);

    // hold D-hl CKB-hl ()
    $hold(negedge CKB, negedge D, 1.0, notifier);

    // mpw CKB-lh NS-lh ()
    $width(posedge CKB, 1.0, 0, notifier);

    // mpw CKB-hl NS-hl ()
    $width(negedge CKB, 1.0, 0, notifier);

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HDFCM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:11:16 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HDFCM8N(D, CKB, Q, QB);
  input D, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (1.0, 1.0);

    // arc CKB --> QB
    (negedge CKB => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CKB-hl ()
    $setup(posedge D, negedge CKB, 1.0, notifier);

    // setup D-hl CKB-hl ()
    $setup(negedge D, negedge CKB, 1.0, notifier);

    // hold D-lh CKB-hl ()
    $hold(negedge CKB, posedge D, 1.0, notifier);

    // hold D-hl CKB-hl ()
    $hold(negedge CKB, negedge D, 1.0, notifier);

    // mpw CKB-lh NS-lh ()
    $width(posedge CKB, 1.0, 0, notifier);

    // mpw CKB-hl NS-hl ()
    $width(negedge CKB, 1.0, 0, notifier);

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HDFCM8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:05:42 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HDFCRSM1N(D, RB, SB, CKB, Q, QB);
  input D, RB, SB, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

    inv_clr0 SMC_I1(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ));

  `ifdef functional // functional //
    dff_p1 SMC_I3(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(RB),
        .preset(SB));

  `else // functional //
    dff_p1 SMC_I3(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(RB), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I5(Q, SMC_IQ);

    buf SMC_I6(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I7(shcheckCKBDhl, RB, SB);

    buf SMC_I8(shcheckCKBRBhl, SB);

    buf SMC_I9(shcheckCKBSBhl, RB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (1.0, 1.0);

    // arc CKB --> QB
    (negedge CKB => ( QB +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl CKB-hl (RB&SB)
    $setup(negedge D &&& (shcheckCKBDhl === 1'b1),
        negedge CKB &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // setup D-lh CKB-hl (RB&SB)
    $setup(posedge D &&& (shcheckCKBDhl === 1'b1),
        negedge CKB &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // setup SB-lh RB-lh ()
    $setup(posedge SB, posedge RB, 1.0, notifier);

    // hold D-hl CKB-hl (RB&SB)
    $hold(negedge CKB &&& (shcheckCKBDhl === 1'b1),
        negedge D &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // hold D-lh CKB-hl (RB&SB)
    $hold(negedge CKB &&& (shcheckCKBDhl === 1'b1),
        posedge D &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // hold SB-lh RB-lh ()
    $hold(posedge RB, posedge SB, 1.0, notifier);

    // recovery RB-lh CKB-hl (SB)
    $recovery(posedge RB &&& (shcheckCKBRBhl === 1'b1),
        negedge CKB &&& (shcheckCKBRBhl === 1'b1), 1.0, notifier);

    // recovery SB-lh CKB-hl (RB)
    $recovery(posedge SB &&& (shcheckCKBSBhl === 1'b1),
        negedge CKB &&& (shcheckCKBSBhl === 1'b1), 1.0, notifier);

    // removal RB-lh CKB-hl (SB)
    $hold(negedge CKB &&& (shcheckCKBRBhl === 1'b1),
        posedge RB &&& (shcheckCKBRBhl === 1'b1), 1.0, notifier);

    // removal SB-lh CKB-hl (RB)
    $hold(negedge CKB &&& (shcheckCKBSBhl === 1'b1),
        posedge SB &&& (shcheckCKBSBhl === 1'b1), 1.0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    // mpw CKB-lh NS-lh ()
    $width(posedge CKB, 1.0, 0, notifier);

    // mpw CKB-hl NS-hl ()
    $width(negedge CKB, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HDFCRSM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:06:30 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HDFCRSM2N(D, RB, SB, CKB, Q, QB);
  input D, RB, SB, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

    inv_clr0 SMC_I1(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ));

  `ifdef functional // functional //
    dff_p1 SMC_I3(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(RB),
        .preset(SB));

  `else // functional //
    dff_p1 SMC_I3(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(RB), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I5(Q, SMC_IQ);

    buf SMC_I6(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I7(shcheckCKBDhl, RB, SB);

    buf SMC_I8(shcheckCKBRBhl, SB);

    buf SMC_I9(shcheckCKBSBhl, RB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (1.0, 1.0);

    // arc CKB --> QB
    (negedge CKB => ( QB +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl CKB-hl (RB&SB)
    $setup(negedge D &&& (shcheckCKBDhl === 1'b1),
        negedge CKB &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // setup D-lh CKB-hl (RB&SB)
    $setup(posedge D &&& (shcheckCKBDhl === 1'b1),
        negedge CKB &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // setup SB-lh RB-lh ()
    $setup(posedge SB, posedge RB, 1.0, notifier);

    // hold D-hl CKB-hl (RB&SB)
    $hold(negedge CKB &&& (shcheckCKBDhl === 1'b1),
        negedge D &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // hold D-lh CKB-hl (RB&SB)
    $hold(negedge CKB &&& (shcheckCKBDhl === 1'b1),
        posedge D &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // hold SB-lh RB-lh ()
    $hold(posedge RB, posedge SB, 1.0, notifier);

    // recovery RB-lh CKB-hl (SB)
    $recovery(posedge RB &&& (shcheckCKBRBhl === 1'b1),
        negedge CKB &&& (shcheckCKBRBhl === 1'b1), 1.0, notifier);

    // recovery SB-lh CKB-hl (RB)
    $recovery(posedge SB &&& (shcheckCKBSBhl === 1'b1),
        negedge CKB &&& (shcheckCKBSBhl === 1'b1), 1.0, notifier);

    // removal RB-lh CKB-hl (SB)
    $hold(negedge CKB &&& (shcheckCKBRBhl === 1'b1),
        posedge RB &&& (shcheckCKBRBhl === 1'b1), 1.0, notifier);

    // removal SB-lh CKB-hl (RB)
    $hold(negedge CKB &&& (shcheckCKBSBhl === 1'b1),
        posedge SB &&& (shcheckCKBSBhl === 1'b1), 1.0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    // mpw CKB-lh NS-lh ()
    $width(posedge CKB, 1.0, 0, notifier);

    // mpw CKB-hl NS-hl ()
    $width(negedge CKB, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HDFCRSM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:12:48 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HDFCRSM4N(D, RB, SB, CKB, Q, QB);
  input D, RB, SB, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

    inv_clr0 SMC_I1(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ));

  `ifdef functional // functional //
    dff_p1 SMC_I3(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(RB),
        .preset(SB));

  `else // functional //
    dff_p1 SMC_I3(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(RB), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I5(Q, SMC_IQ);

    buf SMC_I6(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I7(shcheckCKBDhl, RB, SB);

    buf SMC_I8(shcheckCKBRBhl, SB);

    buf SMC_I9(shcheckCKBSBhl, RB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (1.0, 1.0);

    // arc CKB --> QB
    (negedge CKB => ( QB +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl CKB-hl (RB&SB)
    $setup(negedge D &&& (shcheckCKBDhl === 1'b1),
        negedge CKB &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // setup D-lh CKB-hl (RB&SB)
    $setup(posedge D &&& (shcheckCKBDhl === 1'b1),
        negedge CKB &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // setup SB-lh RB-lh ()
    $setup(posedge SB, posedge RB, 1.0, notifier);

    // hold D-hl CKB-hl (RB&SB)
    $hold(negedge CKB &&& (shcheckCKBDhl === 1'b1),
        negedge D &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // hold D-lh CKB-hl (RB&SB)
    $hold(negedge CKB &&& (shcheckCKBDhl === 1'b1),
        posedge D &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // hold SB-lh RB-lh ()
    $hold(posedge RB, posedge SB, 1.0, notifier);

    // recovery RB-lh CKB-hl (SB)
    $recovery(posedge RB &&& (shcheckCKBRBhl === 1'b1),
        negedge CKB &&& (shcheckCKBRBhl === 1'b1), 1.0, notifier);

    // recovery SB-lh CKB-hl (RB)
    $recovery(posedge SB &&& (shcheckCKBSBhl === 1'b1),
        negedge CKB &&& (shcheckCKBSBhl === 1'b1), 1.0, notifier);

    // removal RB-lh CKB-hl (SB)
    $hold(negedge CKB &&& (shcheckCKBRBhl === 1'b1),
        posedge RB &&& (shcheckCKBRBhl === 1'b1), 1.0, notifier);

    // removal SB-lh CKB-hl (RB)
    $hold(negedge CKB &&& (shcheckCKBSBhl === 1'b1),
        posedge SB &&& (shcheckCKBSBhl === 1'b1), 1.0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    // mpw CKB-lh NS-lh ()
    $width(posedge CKB, 1.0, 0, notifier);

    // mpw CKB-hl NS-hl ()
    $width(negedge CKB, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HDFCRSM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:10:21 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HDFCRSM8N(D, RB, SB, CKB, Q, QB);
  input D, RB, SB, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

    inv_clr0 SMC_I1(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ));

  `ifdef functional // functional //
    dff_p1 SMC_I3(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(RB),
        .preset(SB));

  `else // functional //
    dff_p1 SMC_I3(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(RB), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I5(Q, SMC_IQ);

    buf SMC_I6(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I7(shcheckCKBDhl, RB, SB);

    buf SMC_I8(shcheckCKBRBhl, SB);

    buf SMC_I9(shcheckCKBSBhl, RB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (1.0, 1.0);

    // arc CKB --> QB
    (negedge CKB => ( QB +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl CKB-hl (RB&SB)
    $setup(negedge D &&& (shcheckCKBDhl === 1'b1),
        negedge CKB &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // setup D-lh CKB-hl (RB&SB)
    $setup(posedge D &&& (shcheckCKBDhl === 1'b1),
        negedge CKB &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // setup SB-lh RB-lh ()
    $setup(posedge SB, posedge RB, 1.0, notifier);

    // hold D-hl CKB-hl (RB&SB)
    $hold(negedge CKB &&& (shcheckCKBDhl === 1'b1),
        negedge D &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // hold D-lh CKB-hl (RB&SB)
    $hold(negedge CKB &&& (shcheckCKBDhl === 1'b1),
        posedge D &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // hold SB-lh RB-lh ()
    $hold(posedge RB, posedge SB, 1.0, notifier);

    // recovery RB-lh CKB-hl (SB)
    $recovery(posedge RB &&& (shcheckCKBRBhl === 1'b1),
        negedge CKB &&& (shcheckCKBRBhl === 1'b1), 1.0, notifier);

    // recovery SB-lh CKB-hl (RB)
    $recovery(posedge SB &&& (shcheckCKBSBhl === 1'b1),
        negedge CKB &&& (shcheckCKBSBhl === 1'b1), 1.0, notifier);

    // removal RB-lh CKB-hl (SB)
    $hold(negedge CKB &&& (shcheckCKBRBhl === 1'b1),
        posedge RB &&& (shcheckCKBRBhl === 1'b1), 1.0, notifier);

    // removal SB-lh CKB-hl (RB)
    $hold(negedge CKB &&& (shcheckCKBSBhl === 1'b1),
        posedge SB &&& (shcheckCKBSBhl === 1'b1), 1.0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    // mpw CKB-lh NS-lh ()
    $width(posedge CKB, 1.0, 0, notifier);

    // mpw CKB-hl NS-hl ()
    $width(negedge CKB, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HDFCRSM8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:11:51 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HDFEQM1N(D, E, CK, Q);
  input D, E, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, D, SMC_IQ, E);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I4(shcheckCKDlh, E);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: E )) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // setup D-hl CK-lh (E)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (E)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // hold D-hl CK-lh (E)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (E)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HDFEQM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:10:54 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HDFEQM2N(D, E, CK, Q);
  input D, E, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, D, SMC_IQ, E);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I4(shcheckCKDlh, E);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: E )) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // setup D-hl CK-lh (E)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (E)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // hold D-hl CK-lh (E)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (E)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HDFEQM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:08:51 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HDFEQM4N(D, E, CK, Q);
  input D, E, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, D, SMC_IQ, E);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I4(shcheckCKDlh, E);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: E )) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // setup D-hl CK-lh (E)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (E)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // hold D-hl CK-lh (E)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (E)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HDFEQM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:06:40 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HDFEQM8N(D, E, CK, Q);
  input D, E, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, D, SMC_IQ, E);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I4(shcheckCKDlh, E);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: E )) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // setup D-hl CK-lh (E)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (E)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // hold D-hl CK-lh (E)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (E)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HDFEQM8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:11:22 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HDFM1N(D, CK, Q, QB);
  input D, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh ()
    $setup(posedge D, posedge CK, 1.0, notifier);

    // setup D-hl CK-lh ()
    $setup(negedge D, posedge CK, 1.0, notifier);

    // hold D-lh CK-lh ()
    $hold(posedge CK, posedge D, 1.0, notifier);

    // hold D-hl CK-lh ()
    $hold(posedge CK, negedge D, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HDFM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:08:09 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HDFM2N(D, CK, Q, QB);
  input D, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh ()
    $setup(posedge D, posedge CK, 1.0, notifier);

    // setup D-hl CK-lh ()
    $setup(negedge D, posedge CK, 1.0, notifier);

    // hold D-lh CK-lh ()
    $hold(posedge CK, posedge D, 1.0, notifier);

    // hold D-hl CK-lh ()
    $hold(posedge CK, negedge D, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HDFM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:12:50 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HDFM4N(D, CK, Q, QB);
  input D, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh ()
    $setup(posedge D, posedge CK, 1.0, notifier);

    // setup D-hl CK-lh ()
    $setup(negedge D, posedge CK, 1.0, notifier);

    // hold D-lh CK-lh ()
    $hold(posedge CK, posedge D, 1.0, notifier);

    // hold D-hl CK-lh ()
    $hold(posedge CK, negedge D, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HDFM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:10:35 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HDFM8N(D, CK, Q, QB);
  input D, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh ()
    $setup(posedge D, posedge CK, 1.0, notifier);

    // setup D-hl CK-lh ()
    $setup(negedge D, posedge CK, 1.0, notifier);

    // hold D-lh CK-lh ()
    $hold(posedge CK, posedge D, 1.0, notifier);

    // hold D-hl CK-lh ()
    $hold(posedge CK, negedge D, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HDFM8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:11:59 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HDFMQM1N(D1, D2, S, CK, Q);
  input D1, D2, S, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, D2, D1, S);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(shcheckCKD1lh, S);

    buf SMC_I5(shcheckCKD2lh, S);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D1 )) = (1.0, 1.0);



    // setup S-lh CK-lh ()
    $setup(posedge S, posedge CK, 1.0, notifier);

    // setup S-hl CK-lh ()
    $setup(negedge S, posedge CK, 1.0, notifier);

    // setup D2-lh CK-lh (S)
    $setup(posedge D2 &&& (shcheckCKD2lh === 1'b1),
        posedge CK &&& (shcheckCKD2lh === 1'b1), 1.0, notifier);

    // setup D2-hl CK-lh (S)
    $setup(negedge D2 &&& (shcheckCKD2lh === 1'b1),
        posedge CK &&& (shcheckCKD2lh === 1'b1), 1.0, notifier);

    // setup D1-hl CK-lh (!S)
    $setup(negedge D1 &&& (shcheckCKD1lh === 1'b1),
        posedge CK &&& (shcheckCKD1lh === 1'b1), 1.0, notifier);

    // setup D1-lh CK-lh (!S)
    $setup(posedge D1 &&& (shcheckCKD1lh === 1'b1),
        posedge CK &&& (shcheckCKD1lh === 1'b1), 1.0, notifier);

    // hold S-lh CK-lh ()
    $hold(posedge CK, posedge S, 1.0, notifier);

    // hold S-hl CK-lh ()
    $hold(posedge CK, negedge S, 1.0, notifier);

    // hold D2-lh CK-lh (S)
    $hold(posedge CK &&& (shcheckCKD2lh === 1'b1),
        posedge D2 &&& (shcheckCKD2lh === 1'b1), 1.0, notifier);

    // hold D2-hl CK-lh (S)
    $hold(posedge CK &&& (shcheckCKD2lh === 1'b1),
        negedge D2 &&& (shcheckCKD2lh === 1'b1), 1.0, notifier);

    // hold D1-hl CK-lh (!S)
    $hold(posedge CK &&& (shcheckCKD1lh === 1'b1),
        negedge D1 &&& (shcheckCKD1lh === 1'b1), 1.0, notifier);

    // hold D1-lh CK-lh (!S)
    $hold(posedge CK &&& (shcheckCKD1lh === 1'b1),
        posedge D1 &&& (shcheckCKD1lh === 1'b1), 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HDFMQM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:11:05 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HDFMQM2N(D1, D2, S, CK, Q);
  input D1, D2, S, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, D2, D1, S);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(shcheckCKD1lh, S);

    buf SMC_I5(shcheckCKD2lh, S);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D1 )) = (1.0, 1.0);



    // setup S-lh CK-lh ()
    $setup(posedge S, posedge CK, 1.0, notifier);

    // setup S-hl CK-lh ()
    $setup(negedge S, posedge CK, 1.0, notifier);

    // setup D2-lh CK-lh (S)
    $setup(posedge D2 &&& (shcheckCKD2lh === 1'b1),
        posedge CK &&& (shcheckCKD2lh === 1'b1), 1.0, notifier);

    // setup D2-hl CK-lh (S)
    $setup(negedge D2 &&& (shcheckCKD2lh === 1'b1),
        posedge CK &&& (shcheckCKD2lh === 1'b1), 1.0, notifier);

    // setup D1-hl CK-lh (!S)
    $setup(negedge D1 &&& (shcheckCKD1lh === 1'b1),
        posedge CK &&& (shcheckCKD1lh === 1'b1), 1.0, notifier);

    // setup D1-lh CK-lh (!S)
    $setup(posedge D1 &&& (shcheckCKD1lh === 1'b1),
        posedge CK &&& (shcheckCKD1lh === 1'b1), 1.0, notifier);

    // hold S-lh CK-lh ()
    $hold(posedge CK, posedge S, 1.0, notifier);

    // hold S-hl CK-lh ()
    $hold(posedge CK, negedge S, 1.0, notifier);

    // hold D2-lh CK-lh (S)
    $hold(posedge CK &&& (shcheckCKD2lh === 1'b1),
        posedge D2 &&& (shcheckCKD2lh === 1'b1), 1.0, notifier);

    // hold D2-hl CK-lh (S)
    $hold(posedge CK &&& (shcheckCKD2lh === 1'b1),
        negedge D2 &&& (shcheckCKD2lh === 1'b1), 1.0, notifier);

    // hold D1-hl CK-lh (!S)
    $hold(posedge CK &&& (shcheckCKD1lh === 1'b1),
        negedge D1 &&& (shcheckCKD1lh === 1'b1), 1.0, notifier);

    // hold D1-lh CK-lh (!S)
    $hold(posedge CK &&& (shcheckCKD1lh === 1'b1),
        posedge D1 &&& (shcheckCKD1lh === 1'b1), 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HDFMQM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:06:02 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HDFMQM4N(D1, D2, S, CK, Q);
  input D1, D2, S, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, D2, D1, S);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(shcheckCKD1lh, S);

    buf SMC_I5(shcheckCKD2lh, S);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D1 )) = (1.0, 1.0);



    // setup S-lh CK-lh ()
    $setup(posedge S, posedge CK, 1.0, notifier);

    // setup S-hl CK-lh ()
    $setup(negedge S, posedge CK, 1.0, notifier);

    // setup D2-lh CK-lh (S)
    $setup(posedge D2 &&& (shcheckCKD2lh === 1'b1),
        posedge CK &&& (shcheckCKD2lh === 1'b1), 1.0, notifier);

    // setup D2-hl CK-lh (S)
    $setup(negedge D2 &&& (shcheckCKD2lh === 1'b1),
        posedge CK &&& (shcheckCKD2lh === 1'b1), 1.0, notifier);

    // setup D1-hl CK-lh (!S)
    $setup(negedge D1 &&& (shcheckCKD1lh === 1'b1),
        posedge CK &&& (shcheckCKD1lh === 1'b1), 1.0, notifier);

    // setup D1-lh CK-lh (!S)
    $setup(posedge D1 &&& (shcheckCKD1lh === 1'b1),
        posedge CK &&& (shcheckCKD1lh === 1'b1), 1.0, notifier);

    // hold S-lh CK-lh ()
    $hold(posedge CK, posedge S, 1.0, notifier);

    // hold S-hl CK-lh ()
    $hold(posedge CK, negedge S, 1.0, notifier);

    // hold D2-lh CK-lh (S)
    $hold(posedge CK &&& (shcheckCKD2lh === 1'b1),
        posedge D2 &&& (shcheckCKD2lh === 1'b1), 1.0, notifier);

    // hold D2-hl CK-lh (S)
    $hold(posedge CK &&& (shcheckCKD2lh === 1'b1),
        negedge D2 &&& (shcheckCKD2lh === 1'b1), 1.0, notifier);

    // hold D1-hl CK-lh (!S)
    $hold(posedge CK &&& (shcheckCKD1lh === 1'b1),
        negedge D1 &&& (shcheckCKD1lh === 1'b1), 1.0, notifier);

    // hold D1-lh CK-lh (!S)
    $hold(posedge CK &&& (shcheckCKD1lh === 1'b1),
        posedge D1 &&& (shcheckCKD1lh === 1'b1), 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HDFMQM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:05:57 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HDFMQM8N(D1, D2, S, CK, Q);
  input D1, D2, S, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, D2, D1, S);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(shcheckCKD1lh, S);

    buf SMC_I5(shcheckCKD2lh, S);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D1 )) = (1.0, 1.0);



    // setup S-lh CK-lh ()
    $setup(posedge S, posedge CK, 1.0, notifier);

    // setup S-hl CK-lh ()
    $setup(negedge S, posedge CK, 1.0, notifier);

    // setup D2-lh CK-lh (S)
    $setup(posedge D2 &&& (shcheckCKD2lh === 1'b1),
        posedge CK &&& (shcheckCKD2lh === 1'b1), 1.0, notifier);

    // setup D2-hl CK-lh (S)
    $setup(negedge D2 &&& (shcheckCKD2lh === 1'b1),
        posedge CK &&& (shcheckCKD2lh === 1'b1), 1.0, notifier);

    // setup D1-hl CK-lh (!S)
    $setup(negedge D1 &&& (shcheckCKD1lh === 1'b1),
        posedge CK &&& (shcheckCKD1lh === 1'b1), 1.0, notifier);

    // setup D1-lh CK-lh (!S)
    $setup(posedge D1 &&& (shcheckCKD1lh === 1'b1),
        posedge CK &&& (shcheckCKD1lh === 1'b1), 1.0, notifier);

    // hold S-lh CK-lh ()
    $hold(posedge CK, posedge S, 1.0, notifier);

    // hold S-hl CK-lh ()
    $hold(posedge CK, negedge S, 1.0, notifier);

    // hold D2-lh CK-lh (S)
    $hold(posedge CK &&& (shcheckCKD2lh === 1'b1),
        posedge D2 &&& (shcheckCKD2lh === 1'b1), 1.0, notifier);

    // hold D2-hl CK-lh (S)
    $hold(posedge CK &&& (shcheckCKD2lh === 1'b1),
        negedge D2 &&& (shcheckCKD2lh === 1'b1), 1.0, notifier);

    // hold D1-hl CK-lh (!S)
    $hold(posedge CK &&& (shcheckCKD1lh === 1'b1),
        negedge D1 &&& (shcheckCKD1lh === 1'b1), 1.0, notifier);

    // hold D1-lh CK-lh (!S)
    $hold(posedge CK &&& (shcheckCKD1lh === 1'b1),
        posedge D1 &&& (shcheckCKD1lh === 1'b1), 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HDFMQM8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:06:04 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HDFQM1N(D, CK, Q);
  input D, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh ()
    $setup(negedge D, posedge CK, 1.0, notifier);

    // setup D-lh CK-lh ()
    $setup(posedge D, posedge CK, 1.0, notifier);

    // hold D-hl CK-lh ()
    $hold(posedge CK, negedge D, 1.0, notifier);

    // hold D-lh CK-lh ()
    $hold(posedge CK, posedge D, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HDFQM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:05:58 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HDFQM2N(D, CK, Q);
  input D, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh ()
    $setup(negedge D, posedge CK, 1.0, notifier);

    // setup D-lh CK-lh ()
    $setup(posedge D, posedge CK, 1.0, notifier);

    // hold D-hl CK-lh ()
    $hold(posedge CK, negedge D, 1.0, notifier);

    // hold D-lh CK-lh ()
    $hold(posedge CK, posedge D, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HDFQM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:08:20 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HDFQM4N(D, CK, Q);
  input D, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh ()
    $setup(negedge D, posedge CK, 1.0, notifier);

    // setup D-lh CK-lh ()
    $setup(posedge D, posedge CK, 1.0, notifier);

    // hold D-hl CK-lh ()
    $hold(posedge CK, negedge D, 1.0, notifier);

    // hold D-lh CK-lh ()
    $hold(posedge CK, posedge D, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HDFQM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:13:01 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HDFQM8N(D, CK, Q);
  input D, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh ()
    $setup(negedge D, posedge CK, 1.0, notifier);

    // setup D-lh CK-lh ()
    $setup(posedge D, posedge CK, 1.0, notifier);

    // hold D-hl CK-lh ()
    $hold(posedge CK, negedge D, 1.0, notifier);

    // hold D-lh CK-lh ()
    $hold(posedge CK, posedge D, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HDFQM8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:08:56 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HDFQRM1N(D, RB, CK, Q);
  input D, RB, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckCKDlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (RB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (RB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 1.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HDFQRM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:11:28 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HDFQRM2N(D, RB, CK, Q);
  input D, RB, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckCKDlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (RB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (RB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 1.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HDFQRM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:08:21 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HDFQRM4N(D, RB, CK, Q);
  input D, RB, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckCKDlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (RB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (RB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 1.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HDFQRM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:13:01 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HDFQRM8N(D, RB, CK, Q);
  input D, RB, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckCKDlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (RB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (RB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 1.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HDFQRM8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:10:44 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HDFQRSM1N(D, RB, SB, CK, Q);
  input D, RB, SB, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //
    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(SB));

  `else // functional //
    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I3(shcheckCKDlh, RB, SB);

    buf SMC_I4(shcheckCKRBlh, SB);

    buf SMC_I5(shcheckCKSBlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);



    // setup SB-lh RB-lh ()
    $setup(posedge SB, posedge RB, 1.0, notifier);

    // setup D-lh CK-lh (RB&SB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (RB&SB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SB-lh RB-lh ()
    $hold(posedge RB, posedge SB, 1.0, notifier);

    // hold D-lh CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh (RB)
    $recovery(posedge SB &&& (shcheckCKSBlh === 1'b1),
        posedge CK &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh (SB)
    $recovery(posedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // removal SB-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSBlh === 1'b1),
        posedge SB &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // removal RB-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        posedge RB &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HDFQRSM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:11:12 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HDFQRSM2N(D, RB, SB, CK, Q);
  input D, RB, SB, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //
    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(SB));

  `else // functional //
    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I3(shcheckCKDlh, RB, SB);

    buf SMC_I4(shcheckCKRBlh, SB);

    buf SMC_I5(shcheckCKSBlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);



    // setup SB-lh RB-lh ()
    $setup(posedge SB, posedge RB, 1.0, notifier);

    // setup D-lh CK-lh (RB&SB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (RB&SB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SB-lh RB-lh ()
    $hold(posedge RB, posedge SB, 1.0, notifier);

    // hold D-lh CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh (RB)
    $recovery(posedge SB &&& (shcheckCKSBlh === 1'b1),
        posedge CK &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh (SB)
    $recovery(posedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // removal SB-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSBlh === 1'b1),
        posedge SB &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // removal RB-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        posedge RB &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HDFQRSM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:06:53 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HDFQRSM4N(D, RB, SB, CK, Q);
  input D, RB, SB, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //
    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(SB));

  `else // functional //
    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I3(shcheckCKDlh, RB, SB);

    buf SMC_I4(shcheckCKRBlh, SB);

    buf SMC_I5(shcheckCKSBlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);



    // setup SB-lh RB-lh ()
    $setup(posedge SB, posedge RB, 1.0, notifier);

    // setup D-lh CK-lh (RB&SB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (RB&SB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SB-lh RB-lh ()
    $hold(posedge RB, posedge SB, 1.0, notifier);

    // hold D-lh CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh (RB)
    $recovery(posedge SB &&& (shcheckCKSBlh === 1'b1),
        posedge CK &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh (SB)
    $recovery(posedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // removal SB-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSBlh === 1'b1),
        posedge SB &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // removal RB-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        posedge RB &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HDFQRSM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:09:12 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HDFQRSM8N(D, RB, SB, CK, Q);
  input D, RB, SB, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //
    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(SB));

  `else // functional //
    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I3(shcheckCKDlh, RB, SB);

    buf SMC_I4(shcheckCKRBlh, SB);

    buf SMC_I5(shcheckCKSBlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);



    // setup SB-lh RB-lh ()
    $setup(posedge SB, posedge RB, 1.0, notifier);

    // setup D-lh CK-lh (RB&SB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (RB&SB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SB-lh RB-lh ()
    $hold(posedge RB, posedge SB, 1.0, notifier);

    // hold D-lh CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh (RB)
    $recovery(posedge SB &&& (shcheckCKSBlh === 1'b1),
        posedge CK &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh (SB)
    $recovery(posedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // removal SB-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSBlh === 1'b1),
        posedge SB &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // removal RB-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        posedge RB &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HDFQRSM8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:11:42 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HDFQSM1N(D, SB, CK, Q);
  input D, SB, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //
    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(SB));

  `else // functional //
    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckCKDlh, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (SB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (SB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 1.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HDFQSM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:08:37 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HDFQSM2N(D, SB, CK, Q);
  input D, SB, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //
    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(SB));

  `else // functional //
    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckCKDlh, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (SB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (SB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 1.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HDFQSM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:06:09 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HDFQSM4N(D, SB, CK, Q);
  input D, SB, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //
    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(SB));

  `else // functional //
    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckCKDlh, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (SB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (SB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 1.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HDFQSM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:13:17 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HDFQSM8N(D, SB, CK, Q);
  input D, SB, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //
    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(SB));

  `else // functional //
    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckCKDlh, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (SB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (SB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 1.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HDFQSM8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:12:13 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HSDFCM1N(D, SD, SE, CKB, Q, QB);
  input D, SD, SE, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

    not SMC_I1(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I2(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I5(Q, SMC_IQ);

    buf SMC_I6(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I7(shcheckCKBDhl, SE);

    buf SMC_I8(shcheckCKBSDhl, SE);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (1.0, 1.0);

    // arc CKB --> QB
    (negedge CKB => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CKB-hl (!SE)
    $setup(posedge D &&& (shcheckCKBDhl === 1'b1),
        negedge CKB &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // setup D-hl CKB-hl (!SE)
    $setup(negedge D &&& (shcheckCKBDhl === 1'b1),
        negedge CKB &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // setup SE-lh CKB-hl ()
    $setup(posedge SE, negedge CKB, 1.0, notifier);

    // setup SE-hl CKB-hl ()
    $setup(negedge SE, negedge CKB, 1.0, notifier);

    // setup SD-lh CKB-hl (SE)
    $setup(posedge SD &&& (shcheckCKBSDhl === 1'b1),
        negedge CKB &&& (shcheckCKBSDhl === 1'b1), 1.0, notifier);

    // setup SD-hl CKB-hl (SE)
    $setup(negedge SD &&& (shcheckCKBSDhl === 1'b1),
        negedge CKB &&& (shcheckCKBSDhl === 1'b1), 1.0, notifier);

    // hold D-lh CKB-hl (!SE)
    $hold(negedge CKB &&& (shcheckCKBDhl === 1'b1),
        posedge D &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // hold D-hl CKB-hl (!SE)
    $hold(negedge CKB &&& (shcheckCKBDhl === 1'b1),
        negedge D &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // hold SE-lh CKB-hl ()
    $hold(negedge CKB, posedge SE, 1.0, notifier);

    // hold SE-hl CKB-hl ()
    $hold(negedge CKB, negedge SE, 1.0, notifier);

    // hold SD-lh CKB-hl (SE)
    $hold(negedge CKB &&& (shcheckCKBSDhl === 1'b1),
        posedge SD &&& (shcheckCKBSDhl === 1'b1), 1.0, notifier);

    // hold SD-hl CKB-hl (SE)
    $hold(negedge CKB &&& (shcheckCKBSDhl === 1'b1),
        negedge SD &&& (shcheckCKBSDhl === 1'b1), 1.0, notifier);

    // mpw CKB-lh NS-lh ()
    $width(posedge CKB, 1.0, 0, notifier);

    // mpw CKB-hl NS-hl ()
    $width(negedge CKB, 1.0, 0, notifier);

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HSDFCM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:06:12 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HSDFCM2N(D, SD, SE, CKB, Q, QB);
  input D, SD, SE, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

    not SMC_I1(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I2(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I5(Q, SMC_IQ);

    buf SMC_I6(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I7(shcheckCKBDhl, SE);

    buf SMC_I8(shcheckCKBSDhl, SE);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (1.0, 1.0);

    // arc CKB --> QB
    (negedge CKB => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CKB-hl (!SE)
    $setup(posedge D &&& (shcheckCKBDhl === 1'b1),
        negedge CKB &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // setup D-hl CKB-hl (!SE)
    $setup(negedge D &&& (shcheckCKBDhl === 1'b1),
        negedge CKB &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // setup SE-lh CKB-hl ()
    $setup(posedge SE, negedge CKB, 1.0, notifier);

    // setup SE-hl CKB-hl ()
    $setup(negedge SE, negedge CKB, 1.0, notifier);

    // setup SD-lh CKB-hl (SE)
    $setup(posedge SD &&& (shcheckCKBSDhl === 1'b1),
        negedge CKB &&& (shcheckCKBSDhl === 1'b1), 1.0, notifier);

    // setup SD-hl CKB-hl (SE)
    $setup(negedge SD &&& (shcheckCKBSDhl === 1'b1),
        negedge CKB &&& (shcheckCKBSDhl === 1'b1), 1.0, notifier);

    // hold D-lh CKB-hl (!SE)
    $hold(negedge CKB &&& (shcheckCKBDhl === 1'b1),
        posedge D &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // hold D-hl CKB-hl (!SE)
    $hold(negedge CKB &&& (shcheckCKBDhl === 1'b1),
        negedge D &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // hold SE-lh CKB-hl ()
    $hold(negedge CKB, posedge SE, 1.0, notifier);

    // hold SE-hl CKB-hl ()
    $hold(negedge CKB, negedge SE, 1.0, notifier);

    // hold SD-lh CKB-hl (SE)
    $hold(negedge CKB &&& (shcheckCKBSDhl === 1'b1),
        posedge SD &&& (shcheckCKBSDhl === 1'b1), 1.0, notifier);

    // hold SD-hl CKB-hl (SE)
    $hold(negedge CKB &&& (shcheckCKBSDhl === 1'b1),
        negedge SD &&& (shcheckCKBSDhl === 1'b1), 1.0, notifier);

    // mpw CKB-lh NS-lh ()
    $width(posedge CKB, 1.0, 0, notifier);

    // mpw CKB-hl NS-hl ()
    $width(negedge CKB, 1.0, 0, notifier);

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HSDFCM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:06:12 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HSDFCM4N(D, SD, SE, CKB, Q, QB);
  input D, SD, SE, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

    not SMC_I1(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I2(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I5(Q, SMC_IQ);

    buf SMC_I6(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I7(shcheckCKBDhl, SE);

    buf SMC_I8(shcheckCKBSDhl, SE);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (1.0, 1.0);

    // arc CKB --> QB
    (negedge CKB => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CKB-hl (!SE)
    $setup(posedge D &&& (shcheckCKBDhl === 1'b1),
        negedge CKB &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // setup D-hl CKB-hl (!SE)
    $setup(negedge D &&& (shcheckCKBDhl === 1'b1),
        negedge CKB &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // setup SE-lh CKB-hl ()
    $setup(posedge SE, negedge CKB, 1.0, notifier);

    // setup SE-hl CKB-hl ()
    $setup(negedge SE, negedge CKB, 1.0, notifier);

    // setup SD-lh CKB-hl (SE)
    $setup(posedge SD &&& (shcheckCKBSDhl === 1'b1),
        negedge CKB &&& (shcheckCKBSDhl === 1'b1), 1.0, notifier);

    // setup SD-hl CKB-hl (SE)
    $setup(negedge SD &&& (shcheckCKBSDhl === 1'b1),
        negedge CKB &&& (shcheckCKBSDhl === 1'b1), 1.0, notifier);

    // hold D-lh CKB-hl (!SE)
    $hold(negedge CKB &&& (shcheckCKBDhl === 1'b1),
        posedge D &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // hold D-hl CKB-hl (!SE)
    $hold(negedge CKB &&& (shcheckCKBDhl === 1'b1),
        negedge D &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // hold SE-lh CKB-hl ()
    $hold(negedge CKB, posedge SE, 1.0, notifier);

    // hold SE-hl CKB-hl ()
    $hold(negedge CKB, negedge SE, 1.0, notifier);

    // hold SD-lh CKB-hl (SE)
    $hold(negedge CKB &&& (shcheckCKBSDhl === 1'b1),
        posedge SD &&& (shcheckCKBSDhl === 1'b1), 1.0, notifier);

    // hold SD-hl CKB-hl (SE)
    $hold(negedge CKB &&& (shcheckCKBSDhl === 1'b1),
        negedge SD &&& (shcheckCKBSDhl === 1'b1), 1.0, notifier);

    // mpw CKB-lh NS-lh ()
    $width(posedge CKB, 1.0, 0, notifier);

    // mpw CKB-hl NS-hl ()
    $width(negedge CKB, 1.0, 0, notifier);

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HSDFCM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:11:44 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HSDFCM8N(D, SD, SE, CKB, Q, QB);
  input D, SD, SE, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

    not SMC_I1(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I2(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I5(Q, SMC_IQ);

    buf SMC_I6(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I7(shcheckCKBDhl, SE);

    buf SMC_I8(shcheckCKBSDhl, SE);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (1.0, 1.0);

    // arc CKB --> QB
    (negedge CKB => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CKB-hl (!SE)
    $setup(posedge D &&& (shcheckCKBDhl === 1'b1),
        negedge CKB &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // setup D-hl CKB-hl (!SE)
    $setup(negedge D &&& (shcheckCKBDhl === 1'b1),
        negedge CKB &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // setup SE-lh CKB-hl ()
    $setup(posedge SE, negedge CKB, 1.0, notifier);

    // setup SE-hl CKB-hl ()
    $setup(negedge SE, negedge CKB, 1.0, notifier);

    // setup SD-lh CKB-hl (SE)
    $setup(posedge SD &&& (shcheckCKBSDhl === 1'b1),
        negedge CKB &&& (shcheckCKBSDhl === 1'b1), 1.0, notifier);

    // setup SD-hl CKB-hl (SE)
    $setup(negedge SD &&& (shcheckCKBSDhl === 1'b1),
        negedge CKB &&& (shcheckCKBSDhl === 1'b1), 1.0, notifier);

    // hold D-lh CKB-hl (!SE)
    $hold(negedge CKB &&& (shcheckCKBDhl === 1'b1),
        posedge D &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // hold D-hl CKB-hl (!SE)
    $hold(negedge CKB &&& (shcheckCKBDhl === 1'b1),
        negedge D &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // hold SE-lh CKB-hl ()
    $hold(negedge CKB, posedge SE, 1.0, notifier);

    // hold SE-hl CKB-hl ()
    $hold(negedge CKB, negedge SE, 1.0, notifier);

    // hold SD-lh CKB-hl (SE)
    $hold(negedge CKB &&& (shcheckCKBSDhl === 1'b1),
        posedge SD &&& (shcheckCKBSDhl === 1'b1), 1.0, notifier);

    // hold SD-hl CKB-hl (SE)
    $hold(negedge CKB &&& (shcheckCKBSDhl === 1'b1),
        negedge SD &&& (shcheckCKBSDhl === 1'b1), 1.0, notifier);

    // mpw CKB-lh NS-lh ()
    $width(posedge CKB, 1.0, 0, notifier);

    // mpw CKB-hl NS-hl ()
    $width(negedge CKB, 1.0, 0, notifier);

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HSDFCM8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:09:16 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HSDFCRSM1N(D, RB, SB, SD, SE, CKB, Q, QB);
  input D, RB, SB, SD, SE, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

    inv_clr0 SMC_I1(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ));
  wire SMC_NS_IN;
    mux21 SMC_I3(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p1 SMC_I4(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN), .clear(RB),
        .preset(SB));

  `else // functional //
    dff_p1 SMC_I4(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN), .clear(RB),
        .preset(SB), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I6(Q, SMC_IQ);

    buf SMC_I7(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I8(SE_bar, SE);
    and SMC_I9(shcheckCKBDhl, RB, SB, SE_bar);

    buf SMC_I10(shcheckCKBRBhl, SB);

    buf SMC_I11(shcheckCKBSBhl, RB);

    and SMC_I12(shcheckCKBSDhl, RB, SB, SE);

    and SMC_I13(shcheckCKBSEhl, RB, SB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (1.0, 1.0);

    // arc CKB --> QB
    (negedge CKB => ( QB +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CKB-hl (RB&SB&!SE)
    $setup(posedge D &&& (shcheckCKBDhl === 1'b1),
        negedge CKB &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // setup D-hl CKB-hl (RB&SB&!SE)
    $setup(negedge D &&& (shcheckCKBDhl === 1'b1),
        negedge CKB &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // setup SB-lh RB-lh ()
    $setup(posedge SB, posedge RB, 1.0, notifier);

    // setup SE-hl CKB-hl (RB&SB)
    $setup(negedge SE &&& (shcheckCKBSEhl === 1'b1),
        negedge CKB &&& (shcheckCKBSEhl === 1'b1), 1.0, notifier);

    // setup SE-lh CKB-hl (RB&SB)
    $setup(posedge SE &&& (shcheckCKBSEhl === 1'b1),
        negedge CKB &&& (shcheckCKBSEhl === 1'b1), 1.0, notifier);

    // setup SD-hl CKB-hl (RB&SB&SE)
    $setup(negedge SD &&& (shcheckCKBSDhl === 1'b1),
        negedge CKB &&& (shcheckCKBSDhl === 1'b1), 1.0, notifier);

    // setup SD-lh CKB-hl (RB&SB&SE)
    $setup(posedge SD &&& (shcheckCKBSDhl === 1'b1),
        negedge CKB &&& (shcheckCKBSDhl === 1'b1), 1.0, notifier);

    // hold D-lh CKB-hl (RB&SB&!SE)
    $hold(negedge CKB &&& (shcheckCKBDhl === 1'b1),
        posedge D &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // hold D-hl CKB-hl (RB&SB&!SE)
    $hold(negedge CKB &&& (shcheckCKBDhl === 1'b1),
        negedge D &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // hold SB-lh RB-lh ()
    $hold(posedge RB, posedge SB, 1.0, notifier);

    // hold SE-hl CKB-hl (RB&SB)
    $hold(negedge CKB &&& (shcheckCKBSEhl === 1'b1),
        negedge SE &&& (shcheckCKBSEhl === 1'b1), 1.0, notifier);

    // hold SE-lh CKB-hl (RB&SB)
    $hold(negedge CKB &&& (shcheckCKBSEhl === 1'b1),
        posedge SE &&& (shcheckCKBSEhl === 1'b1), 1.0, notifier);

    // hold SD-hl CKB-hl (RB&SB&SE)
    $hold(negedge CKB &&& (shcheckCKBSDhl === 1'b1),
        negedge SD &&& (shcheckCKBSDhl === 1'b1), 1.0, notifier);

    // hold SD-lh CKB-hl (RB&SB&SE)
    $hold(negedge CKB &&& (shcheckCKBSDhl === 1'b1),
        posedge SD &&& (shcheckCKBSDhl === 1'b1), 1.0, notifier);

    // recovery RB-lh CKB-hl (SB)
    $recovery(posedge RB &&& (shcheckCKBRBhl === 1'b1),
        negedge CKB &&& (shcheckCKBRBhl === 1'b1), 1.0, notifier);

    // recovery SB-lh CKB-hl (RB)
    $recovery(posedge SB &&& (shcheckCKBSBhl === 1'b1),
        negedge CKB &&& (shcheckCKBSBhl === 1'b1), 1.0, notifier);

    // removal RB-lh CKB-hl (SB)
    $hold(negedge CKB &&& (shcheckCKBRBhl === 1'b1),
        posedge RB &&& (shcheckCKBRBhl === 1'b1), 1.0, notifier);

    // removal SB-lh CKB-hl (RB)
    $hold(negedge CKB &&& (shcheckCKBSBhl === 1'b1),
        posedge SB &&& (shcheckCKBSBhl === 1'b1), 1.0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    // mpw CKB-lh NS-lh ()
    $width(posedge CKB, 1.0, 0, notifier);

    // mpw CKB-hl NS-hl ()
    $width(negedge CKB, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HSDFCRSM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:06:58 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HSDFCRSM2N(D, RB, SB, SD, SE, CKB, Q, QB);
  input D, RB, SB, SD, SE, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

    inv_clr0 SMC_I1(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ));
  wire SMC_NS_IN;
    mux21 SMC_I3(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p1 SMC_I4(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN), .clear(RB),
        .preset(SB));

  `else // functional //
    dff_p1 SMC_I4(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN), .clear(RB),
        .preset(SB), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I6(Q, SMC_IQ);

    buf SMC_I7(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I8(SE_bar, SE);
    and SMC_I9(shcheckCKBDhl, RB, SB, SE_bar);

    buf SMC_I10(shcheckCKBRBhl, SB);

    buf SMC_I11(shcheckCKBSBhl, RB);

    and SMC_I12(shcheckCKBSDhl, RB, SB, SE);

    and SMC_I13(shcheckCKBSEhl, RB, SB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (1.0, 1.0);

    // arc CKB --> QB
    (negedge CKB => ( QB +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CKB-hl (RB&SB&!SE)
    $setup(posedge D &&& (shcheckCKBDhl === 1'b1),
        negedge CKB &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // setup D-hl CKB-hl (RB&SB&!SE)
    $setup(negedge D &&& (shcheckCKBDhl === 1'b1),
        negedge CKB &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // setup SB-lh RB-lh ()
    $setup(posedge SB, posedge RB, 1.0, notifier);

    // setup SE-hl CKB-hl (RB&SB)
    $setup(negedge SE &&& (shcheckCKBSEhl === 1'b1),
        negedge CKB &&& (shcheckCKBSEhl === 1'b1), 1.0, notifier);

    // setup SE-lh CKB-hl (RB&SB)
    $setup(posedge SE &&& (shcheckCKBSEhl === 1'b1),
        negedge CKB &&& (shcheckCKBSEhl === 1'b1), 1.0, notifier);

    // setup SD-hl CKB-hl (RB&SB&SE)
    $setup(negedge SD &&& (shcheckCKBSDhl === 1'b1),
        negedge CKB &&& (shcheckCKBSDhl === 1'b1), 1.0, notifier);

    // setup SD-lh CKB-hl (RB&SB&SE)
    $setup(posedge SD &&& (shcheckCKBSDhl === 1'b1),
        negedge CKB &&& (shcheckCKBSDhl === 1'b1), 1.0, notifier);

    // hold D-lh CKB-hl (RB&SB&!SE)
    $hold(negedge CKB &&& (shcheckCKBDhl === 1'b1),
        posedge D &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // hold D-hl CKB-hl (RB&SB&!SE)
    $hold(negedge CKB &&& (shcheckCKBDhl === 1'b1),
        negedge D &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // hold SB-lh RB-lh ()
    $hold(posedge RB, posedge SB, 1.0, notifier);

    // hold SE-hl CKB-hl (RB&SB)
    $hold(negedge CKB &&& (shcheckCKBSEhl === 1'b1),
        negedge SE &&& (shcheckCKBSEhl === 1'b1), 1.0, notifier);

    // hold SE-lh CKB-hl (RB&SB)
    $hold(negedge CKB &&& (shcheckCKBSEhl === 1'b1),
        posedge SE &&& (shcheckCKBSEhl === 1'b1), 1.0, notifier);

    // hold SD-hl CKB-hl (RB&SB&SE)
    $hold(negedge CKB &&& (shcheckCKBSDhl === 1'b1),
        negedge SD &&& (shcheckCKBSDhl === 1'b1), 1.0, notifier);

    // hold SD-lh CKB-hl (RB&SB&SE)
    $hold(negedge CKB &&& (shcheckCKBSDhl === 1'b1),
        posedge SD &&& (shcheckCKBSDhl === 1'b1), 1.0, notifier);

    // recovery RB-lh CKB-hl (SB)
    $recovery(posedge RB &&& (shcheckCKBRBhl === 1'b1),
        negedge CKB &&& (shcheckCKBRBhl === 1'b1), 1.0, notifier);

    // recovery SB-lh CKB-hl (RB)
    $recovery(posedge SB &&& (shcheckCKBSBhl === 1'b1),
        negedge CKB &&& (shcheckCKBSBhl === 1'b1), 1.0, notifier);

    // removal RB-lh CKB-hl (SB)
    $hold(negedge CKB &&& (shcheckCKBRBhl === 1'b1),
        posedge RB &&& (shcheckCKBRBhl === 1'b1), 1.0, notifier);

    // removal SB-lh CKB-hl (RB)
    $hold(negedge CKB &&& (shcheckCKBSBhl === 1'b1),
        posedge SB &&& (shcheckCKBSBhl === 1'b1), 1.0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    // mpw CKB-lh NS-lh ()
    $width(posedge CKB, 1.0, 0, notifier);

    // mpw CKB-hl NS-hl ()
    $width(negedge CKB, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HSDFCRSM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:09:00 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HSDFCRSM4N(D, RB, SB, SD, SE, CKB, Q, QB);
  input D, RB, SB, SD, SE, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

    inv_clr0 SMC_I1(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ));
  wire SMC_NS_IN;
    mux21 SMC_I3(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p1 SMC_I4(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN), .clear(RB),
        .preset(SB));

  `else // functional //
    dff_p1 SMC_I4(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN), .clear(RB),
        .preset(SB), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I6(Q, SMC_IQ);

    buf SMC_I7(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I8(SE_bar, SE);
    and SMC_I9(shcheckCKBDhl, RB, SB, SE_bar);

    buf SMC_I10(shcheckCKBRBhl, SB);

    buf SMC_I11(shcheckCKBSBhl, RB);

    and SMC_I12(shcheckCKBSDhl, RB, SB, SE);

    and SMC_I13(shcheckCKBSEhl, RB, SB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (1.0, 1.0);

    // arc CKB --> QB
    (negedge CKB => ( QB +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CKB-hl (RB&SB&!SE)
    $setup(posedge D &&& (shcheckCKBDhl === 1'b1),
        negedge CKB &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // setup D-hl CKB-hl (RB&SB&!SE)
    $setup(negedge D &&& (shcheckCKBDhl === 1'b1),
        negedge CKB &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // setup SB-lh RB-lh ()
    $setup(posedge SB, posedge RB, 1.0, notifier);

    // setup SE-hl CKB-hl (RB&SB)
    $setup(negedge SE &&& (shcheckCKBSEhl === 1'b1),
        negedge CKB &&& (shcheckCKBSEhl === 1'b1), 1.0, notifier);

    // setup SE-lh CKB-hl (RB&SB)
    $setup(posedge SE &&& (shcheckCKBSEhl === 1'b1),
        negedge CKB &&& (shcheckCKBSEhl === 1'b1), 1.0, notifier);

    // setup SD-hl CKB-hl (RB&SB&SE)
    $setup(negedge SD &&& (shcheckCKBSDhl === 1'b1),
        negedge CKB &&& (shcheckCKBSDhl === 1'b1), 1.0, notifier);

    // setup SD-lh CKB-hl (RB&SB&SE)
    $setup(posedge SD &&& (shcheckCKBSDhl === 1'b1),
        negedge CKB &&& (shcheckCKBSDhl === 1'b1), 1.0, notifier);

    // hold D-lh CKB-hl (RB&SB&!SE)
    $hold(negedge CKB &&& (shcheckCKBDhl === 1'b1),
        posedge D &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // hold D-hl CKB-hl (RB&SB&!SE)
    $hold(negedge CKB &&& (shcheckCKBDhl === 1'b1),
        negedge D &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // hold SB-lh RB-lh ()
    $hold(posedge RB, posedge SB, 1.0, notifier);

    // hold SE-hl CKB-hl (RB&SB)
    $hold(negedge CKB &&& (shcheckCKBSEhl === 1'b1),
        negedge SE &&& (shcheckCKBSEhl === 1'b1), 1.0, notifier);

    // hold SE-lh CKB-hl (RB&SB)
    $hold(negedge CKB &&& (shcheckCKBSEhl === 1'b1),
        posedge SE &&& (shcheckCKBSEhl === 1'b1), 1.0, notifier);

    // hold SD-hl CKB-hl (RB&SB&SE)
    $hold(negedge CKB &&& (shcheckCKBSDhl === 1'b1),
        negedge SD &&& (shcheckCKBSDhl === 1'b1), 1.0, notifier);

    // hold SD-lh CKB-hl (RB&SB&SE)
    $hold(negedge CKB &&& (shcheckCKBSDhl === 1'b1),
        posedge SD &&& (shcheckCKBSDhl === 1'b1), 1.0, notifier);

    // recovery RB-lh CKB-hl (SB)
    $recovery(posedge RB &&& (shcheckCKBRBhl === 1'b1),
        negedge CKB &&& (shcheckCKBRBhl === 1'b1), 1.0, notifier);

    // recovery SB-lh CKB-hl (RB)
    $recovery(posedge SB &&& (shcheckCKBSBhl === 1'b1),
        negedge CKB &&& (shcheckCKBSBhl === 1'b1), 1.0, notifier);

    // removal RB-lh CKB-hl (SB)
    $hold(negedge CKB &&& (shcheckCKBRBhl === 1'b1),
        posedge RB &&& (shcheckCKBRBhl === 1'b1), 1.0, notifier);

    // removal SB-lh CKB-hl (RB)
    $hold(negedge CKB &&& (shcheckCKBSBhl === 1'b1),
        posedge SB &&& (shcheckCKBSBhl === 1'b1), 1.0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    // mpw CKB-lh NS-lh ()
    $width(posedge CKB, 1.0, 0, notifier);

    // mpw CKB-hl NS-hl ()
    $width(negedge CKB, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HSDFCRSM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:11:44 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HSDFCRSM8N(D, RB, SB, SD, SE, CKB, Q, QB);
  input D, RB, SB, SD, SE, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

    inv_clr0 SMC_I1(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ));
  wire SMC_NS_IN;
    mux21 SMC_I3(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p1 SMC_I4(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN), .clear(RB),
        .preset(SB));

  `else // functional //
    dff_p1 SMC_I4(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN), .clear(RB),
        .preset(SB), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I6(Q, SMC_IQ);

    buf SMC_I7(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I8(SE_bar, SE);
    and SMC_I9(shcheckCKBDhl, RB, SB, SE_bar);

    buf SMC_I10(shcheckCKBRBhl, SB);

    buf SMC_I11(shcheckCKBSBhl, RB);

    and SMC_I12(shcheckCKBSDhl, RB, SB, SE);

    and SMC_I13(shcheckCKBSEhl, RB, SB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (1.0, 1.0);

    // arc CKB --> QB
    (negedge CKB => ( QB +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CKB-hl (RB&SB&!SE)
    $setup(posedge D &&& (shcheckCKBDhl === 1'b1),
        negedge CKB &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // setup D-hl CKB-hl (RB&SB&!SE)
    $setup(negedge D &&& (shcheckCKBDhl === 1'b1),
        negedge CKB &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // setup SB-lh RB-lh ()
    $setup(posedge SB, posedge RB, 1.0, notifier);

    // setup SE-hl CKB-hl (RB&SB)
    $setup(negedge SE &&& (shcheckCKBSEhl === 1'b1),
        negedge CKB &&& (shcheckCKBSEhl === 1'b1), 1.0, notifier);

    // setup SE-lh CKB-hl (RB&SB)
    $setup(posedge SE &&& (shcheckCKBSEhl === 1'b1),
        negedge CKB &&& (shcheckCKBSEhl === 1'b1), 1.0, notifier);

    // setup SD-hl CKB-hl (RB&SB&SE)
    $setup(negedge SD &&& (shcheckCKBSDhl === 1'b1),
        negedge CKB &&& (shcheckCKBSDhl === 1'b1), 1.0, notifier);

    // setup SD-lh CKB-hl (RB&SB&SE)
    $setup(posedge SD &&& (shcheckCKBSDhl === 1'b1),
        negedge CKB &&& (shcheckCKBSDhl === 1'b1), 1.0, notifier);

    // hold D-lh CKB-hl (RB&SB&!SE)
    $hold(negedge CKB &&& (shcheckCKBDhl === 1'b1),
        posedge D &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // hold D-hl CKB-hl (RB&SB&!SE)
    $hold(negedge CKB &&& (shcheckCKBDhl === 1'b1),
        negedge D &&& (shcheckCKBDhl === 1'b1), 1.0, notifier);

    // hold SB-lh RB-lh ()
    $hold(posedge RB, posedge SB, 1.0, notifier);

    // hold SE-hl CKB-hl (RB&SB)
    $hold(negedge CKB &&& (shcheckCKBSEhl === 1'b1),
        negedge SE &&& (shcheckCKBSEhl === 1'b1), 1.0, notifier);

    // hold SE-lh CKB-hl (RB&SB)
    $hold(negedge CKB &&& (shcheckCKBSEhl === 1'b1),
        posedge SE &&& (shcheckCKBSEhl === 1'b1), 1.0, notifier);

    // hold SD-hl CKB-hl (RB&SB&SE)
    $hold(negedge CKB &&& (shcheckCKBSDhl === 1'b1),
        negedge SD &&& (shcheckCKBSDhl === 1'b1), 1.0, notifier);

    // hold SD-lh CKB-hl (RB&SB&SE)
    $hold(negedge CKB &&& (shcheckCKBSDhl === 1'b1),
        posedge SD &&& (shcheckCKBSDhl === 1'b1), 1.0, notifier);

    // recovery RB-lh CKB-hl (SB)
    $recovery(posedge RB &&& (shcheckCKBRBhl === 1'b1),
        negedge CKB &&& (shcheckCKBRBhl === 1'b1), 1.0, notifier);

    // recovery SB-lh CKB-hl (RB)
    $recovery(posedge SB &&& (shcheckCKBSBhl === 1'b1),
        negedge CKB &&& (shcheckCKBSBhl === 1'b1), 1.0, notifier);

    // removal RB-lh CKB-hl (SB)
    $hold(negedge CKB &&& (shcheckCKBRBhl === 1'b1),
        posedge RB &&& (shcheckCKBRBhl === 1'b1), 1.0, notifier);

    // removal SB-lh CKB-hl (RB)
    $hold(negedge CKB &&& (shcheckCKBSBhl === 1'b1),
        posedge SB &&& (shcheckCKBSBhl === 1'b1), 1.0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    // mpw CKB-lh NS-lh ()
    $width(posedge CKB, 1.0, 0, notifier);

    // mpw CKB-hl NS-hl ()
    $width(negedge CKB, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HSDFCRSM8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:12:15 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HSDFEQM1N(D, E, SD, SE, CK, Q);
  input D, E, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    HSDFEQM1N_UDP__OUT__ SMC_I0(SMC_NS_IN, D, E, SMC_IQ, SD, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKDlh, E, SE_bar);

    not SMC_I6(shcheckCKElh, SE);

    buf SMC_I7(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);



    // setup E-lh CK-lh (!SE)
    $setup(posedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // setup E-hl CK-lh (!SE)
    $setup(negedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (E&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (E&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold E-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        posedge E &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // hold E-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        negedge E &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (E&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (E&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HSDFEQM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:13:20 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HSDFEQM2N(D, E, SD, SE, CK, Q);
  input D, E, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    HSDFEQM1N_UDP__OUT__ SMC_I0(SMC_NS_IN, D, E, SMC_IQ, SD, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKDlh, E, SE_bar);

    not SMC_I6(shcheckCKElh, SE);

    buf SMC_I7(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);



    // setup E-lh CK-lh (!SE)
    $setup(posedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // setup E-hl CK-lh (!SE)
    $setup(negedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (E&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (E&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold E-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        posedge E &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // hold E-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        negedge E &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (E&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (E&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HSDFEQM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:11:35 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HSDFEQM4N(D, E, SD, SE, CK, Q);
  input D, E, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    HSDFEQM1N_UDP__OUT__ SMC_I0(SMC_NS_IN, D, E, SMC_IQ, SD, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKDlh, E, SE_bar);

    not SMC_I6(shcheckCKElh, SE);

    buf SMC_I7(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);



    // setup E-lh CK-lh (!SE)
    $setup(posedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // setup E-hl CK-lh (!SE)
    $setup(negedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (E&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (E&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold E-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        posedge E &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // hold E-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        negedge E &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (E&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (E&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HSDFEQM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:11:47 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HSDFEQM8N(D, E, SD, SE, CK, Q);
  input D, E, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    HSDFEQM1N_UDP__OUT__ SMC_I0(SMC_NS_IN, D, E, SMC_IQ, SD, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKDlh, E, SE_bar);

    not SMC_I6(shcheckCKElh, SE);

    buf SMC_I7(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);



    // setup E-lh CK-lh (!SE)
    $setup(posedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // setup E-hl CK-lh (!SE)
    $setup(negedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (E&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (E&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold E-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        posedge E &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // hold E-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        negedge E &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (E&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (E&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HSDFEQM8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:07:43 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HSDFM1N(D, SD, SE, CK, Q, QB);
  input D, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(shcheckCKDlh, SE);

    buf SMC_I7(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HSDFM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:10:02 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HSDFM2N(D, SD, SE, CK, Q, QB);
  input D, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(shcheckCKDlh, SE);

    buf SMC_I7(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HSDFM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:09:30 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HSDFM4N(D, SD, SE, CK, Q, QB);
  input D, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(shcheckCKDlh, SE);

    buf SMC_I7(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HSDFM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:12:09 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HSDFM8N(D, SD, SE, CK, Q, QB);
  input D, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(shcheckCKDlh, SE);

    buf SMC_I7(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HSDFM8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:13:07 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HSDFMQM1N(D1, D2, S, SD, SE, CK, Q);
  input D1, D2, S, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    not SMC_I0(SE_bar, SE);
    and SMC_I1(OUT0, D2, S, SE_bar);
    not SMC_I2(S_bar, S);
    and SMC_I3(OUT1, D1, S_bar, SE_bar);
    and SMC_I4(OUT2, SD, SE);
    or SMC_I5(SMC_NS_IN, OUT0, OUT1, OUT2);


  `ifdef functional // functional //
    dff_p0 SMC_I6(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I6(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I8(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I9(shcheckCKD1lh, S_bar, SE_bar);

    and SMC_I10(shcheckCKD2lh, S, SE_bar);

    buf SMC_I11(shcheckCKSDlh, SE);

    not SMC_I12(shcheckCKSlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D1 )) = (1.0, 1.0);



    // setup S-lh CK-lh (!SE)
    $setup(posedge S &&& (shcheckCKSlh === 1'b1),
        posedge CK &&& (shcheckCKSlh === 1'b1), 1.0, notifier);

    // setup S-hl CK-lh (!SE)
    $setup(negedge S &&& (shcheckCKSlh === 1'b1),
        posedge CK &&& (shcheckCKSlh === 1'b1), 1.0, notifier);

    // setup D1-hl CK-lh (!S&!SE)
    $setup(negedge D1 &&& (shcheckCKD1lh === 1'b1),
        posedge CK &&& (shcheckCKD1lh === 1'b1), 1.0, notifier);

    // setup D1-lh CK-lh (!S&!SE)
    $setup(posedge D1 &&& (shcheckCKD1lh === 1'b1),
        posedge CK &&& (shcheckCKD1lh === 1'b1), 1.0, notifier);

    // setup D2-hl CK-lh (S&!SE)
    $setup(negedge D2 &&& (shcheckCKD2lh === 1'b1),
        posedge CK &&& (shcheckCKD2lh === 1'b1), 1.0, notifier);

    // setup D2-lh CK-lh (S&!SE)
    $setup(posedge D2 &&& (shcheckCKD2lh === 1'b1),
        posedge CK &&& (shcheckCKD2lh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold S-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKSlh === 1'b1),
        posedge S &&& (shcheckCKSlh === 1'b1), 1.0, notifier);

    // hold S-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKSlh === 1'b1),
        negedge S &&& (shcheckCKSlh === 1'b1), 1.0, notifier);

    // hold D1-hl CK-lh (!S&!SE)
    $hold(posedge CK &&& (shcheckCKD1lh === 1'b1),
        negedge D1 &&& (shcheckCKD1lh === 1'b1), 1.0, notifier);

    // hold D1-lh CK-lh (!S&!SE)
    $hold(posedge CK &&& (shcheckCKD1lh === 1'b1),
        posedge D1 &&& (shcheckCKD1lh === 1'b1), 1.0, notifier);

    // hold D2-hl CK-lh (S&!SE)
    $hold(posedge CK &&& (shcheckCKD2lh === 1'b1),
        negedge D2 &&& (shcheckCKD2lh === 1'b1), 1.0, notifier);

    // hold D2-lh CK-lh (S&!SE)
    $hold(posedge CK &&& (shcheckCKD2lh === 1'b1),
        posedge D2 &&& (shcheckCKD2lh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HSDFMQM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:11:05 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HSDFMQM2N(D1, D2, S, SD, SE, CK, Q);
  input D1, D2, S, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    not SMC_I0(SE_bar, SE);
    and SMC_I1(OUT0, D2, S, SE_bar);
    not SMC_I2(S_bar, S);
    and SMC_I3(OUT1, D1, S_bar, SE_bar);
    and SMC_I4(OUT2, SD, SE);
    or SMC_I5(SMC_NS_IN, OUT0, OUT1, OUT2);


  `ifdef functional // functional //
    dff_p0 SMC_I6(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I6(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I8(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I9(shcheckCKD1lh, S_bar, SE_bar);

    and SMC_I10(shcheckCKD2lh, S, SE_bar);

    buf SMC_I11(shcheckCKSDlh, SE);

    not SMC_I12(shcheckCKSlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D1 )) = (1.0, 1.0);



    // setup S-lh CK-lh (!SE)
    $setup(posedge S &&& (shcheckCKSlh === 1'b1),
        posedge CK &&& (shcheckCKSlh === 1'b1), 1.0, notifier);

    // setup S-hl CK-lh (!SE)
    $setup(negedge S &&& (shcheckCKSlh === 1'b1),
        posedge CK &&& (shcheckCKSlh === 1'b1), 1.0, notifier);

    // setup D1-hl CK-lh (!S&!SE)
    $setup(negedge D1 &&& (shcheckCKD1lh === 1'b1),
        posedge CK &&& (shcheckCKD1lh === 1'b1), 1.0, notifier);

    // setup D1-lh CK-lh (!S&!SE)
    $setup(posedge D1 &&& (shcheckCKD1lh === 1'b1),
        posedge CK &&& (shcheckCKD1lh === 1'b1), 1.0, notifier);

    // setup D2-hl CK-lh (S&!SE)
    $setup(negedge D2 &&& (shcheckCKD2lh === 1'b1),
        posedge CK &&& (shcheckCKD2lh === 1'b1), 1.0, notifier);

    // setup D2-lh CK-lh (S&!SE)
    $setup(posedge D2 &&& (shcheckCKD2lh === 1'b1),
        posedge CK &&& (shcheckCKD2lh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold S-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKSlh === 1'b1),
        posedge S &&& (shcheckCKSlh === 1'b1), 1.0, notifier);

    // hold S-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKSlh === 1'b1),
        negedge S &&& (shcheckCKSlh === 1'b1), 1.0, notifier);

    // hold D1-hl CK-lh (!S&!SE)
    $hold(posedge CK &&& (shcheckCKD1lh === 1'b1),
        negedge D1 &&& (shcheckCKD1lh === 1'b1), 1.0, notifier);

    // hold D1-lh CK-lh (!S&!SE)
    $hold(posedge CK &&& (shcheckCKD1lh === 1'b1),
        posedge D1 &&& (shcheckCKD1lh === 1'b1), 1.0, notifier);

    // hold D2-hl CK-lh (S&!SE)
    $hold(posedge CK &&& (shcheckCKD2lh === 1'b1),
        negedge D2 &&& (shcheckCKD2lh === 1'b1), 1.0, notifier);

    // hold D2-lh CK-lh (S&!SE)
    $hold(posedge CK &&& (shcheckCKD2lh === 1'b1),
        posedge D2 &&& (shcheckCKD2lh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HSDFMQM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:13:32 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HSDFMQM4N(D1, D2, S, SD, SE, CK, Q);
  input D1, D2, S, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    not SMC_I0(SE_bar, SE);
    and SMC_I1(OUT0, D2, S, SE_bar);
    not SMC_I2(S_bar, S);
    and SMC_I3(OUT1, D1, S_bar, SE_bar);
    and SMC_I4(OUT2, SD, SE);
    or SMC_I5(SMC_NS_IN, OUT0, OUT1, OUT2);


  `ifdef functional // functional //
    dff_p0 SMC_I6(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I6(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I8(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I9(shcheckCKD1lh, S_bar, SE_bar);

    and SMC_I10(shcheckCKD2lh, S, SE_bar);

    buf SMC_I11(shcheckCKSDlh, SE);

    not SMC_I12(shcheckCKSlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D1 )) = (1.0, 1.0);



    // setup S-lh CK-lh (!SE)
    $setup(posedge S &&& (shcheckCKSlh === 1'b1),
        posedge CK &&& (shcheckCKSlh === 1'b1), 1.0, notifier);

    // setup S-hl CK-lh (!SE)
    $setup(negedge S &&& (shcheckCKSlh === 1'b1),
        posedge CK &&& (shcheckCKSlh === 1'b1), 1.0, notifier);

    // setup D1-hl CK-lh (!S&!SE)
    $setup(negedge D1 &&& (shcheckCKD1lh === 1'b1),
        posedge CK &&& (shcheckCKD1lh === 1'b1), 1.0, notifier);

    // setup D1-lh CK-lh (!S&!SE)
    $setup(posedge D1 &&& (shcheckCKD1lh === 1'b1),
        posedge CK &&& (shcheckCKD1lh === 1'b1), 1.0, notifier);

    // setup D2-hl CK-lh (S&!SE)
    $setup(negedge D2 &&& (shcheckCKD2lh === 1'b1),
        posedge CK &&& (shcheckCKD2lh === 1'b1), 1.0, notifier);

    // setup D2-lh CK-lh (S&!SE)
    $setup(posedge D2 &&& (shcheckCKD2lh === 1'b1),
        posedge CK &&& (shcheckCKD2lh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold S-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKSlh === 1'b1),
        posedge S &&& (shcheckCKSlh === 1'b1), 1.0, notifier);

    // hold S-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKSlh === 1'b1),
        negedge S &&& (shcheckCKSlh === 1'b1), 1.0, notifier);

    // hold D1-hl CK-lh (!S&!SE)
    $hold(posedge CK &&& (shcheckCKD1lh === 1'b1),
        negedge D1 &&& (shcheckCKD1lh === 1'b1), 1.0, notifier);

    // hold D1-lh CK-lh (!S&!SE)
    $hold(posedge CK &&& (shcheckCKD1lh === 1'b1),
        posedge D1 &&& (shcheckCKD1lh === 1'b1), 1.0, notifier);

    // hold D2-hl CK-lh (S&!SE)
    $hold(posedge CK &&& (shcheckCKD2lh === 1'b1),
        negedge D2 &&& (shcheckCKD2lh === 1'b1), 1.0, notifier);

    // hold D2-lh CK-lh (S&!SE)
    $hold(posedge CK &&& (shcheckCKD2lh === 1'b1),
        posedge D2 &&& (shcheckCKD2lh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HSDFMQM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:06:27 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HSDFMQM8N(D1, D2, S, SD, SE, CK, Q);
  input D1, D2, S, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    not SMC_I0(SE_bar, SE);
    and SMC_I1(OUT0, D2, S, SE_bar);
    not SMC_I2(S_bar, S);
    and SMC_I3(OUT1, D1, S_bar, SE_bar);
    and SMC_I4(OUT2, SD, SE);
    or SMC_I5(SMC_NS_IN, OUT0, OUT1, OUT2);


  `ifdef functional // functional //
    dff_p0 SMC_I6(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I6(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I8(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I9(shcheckCKD1lh, S_bar, SE_bar);

    and SMC_I10(shcheckCKD2lh, S, SE_bar);

    buf SMC_I11(shcheckCKSDlh, SE);

    not SMC_I12(shcheckCKSlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D1 )) = (1.0, 1.0);



    // setup S-lh CK-lh (!SE)
    $setup(posedge S &&& (shcheckCKSlh === 1'b1),
        posedge CK &&& (shcheckCKSlh === 1'b1), 1.0, notifier);

    // setup S-hl CK-lh (!SE)
    $setup(negedge S &&& (shcheckCKSlh === 1'b1),
        posedge CK &&& (shcheckCKSlh === 1'b1), 1.0, notifier);

    // setup D1-hl CK-lh (!S&!SE)
    $setup(negedge D1 &&& (shcheckCKD1lh === 1'b1),
        posedge CK &&& (shcheckCKD1lh === 1'b1), 1.0, notifier);

    // setup D1-lh CK-lh (!S&!SE)
    $setup(posedge D1 &&& (shcheckCKD1lh === 1'b1),
        posedge CK &&& (shcheckCKD1lh === 1'b1), 1.0, notifier);

    // setup D2-hl CK-lh (S&!SE)
    $setup(negedge D2 &&& (shcheckCKD2lh === 1'b1),
        posedge CK &&& (shcheckCKD2lh === 1'b1), 1.0, notifier);

    // setup D2-lh CK-lh (S&!SE)
    $setup(posedge D2 &&& (shcheckCKD2lh === 1'b1),
        posedge CK &&& (shcheckCKD2lh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold S-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKSlh === 1'b1),
        posedge S &&& (shcheckCKSlh === 1'b1), 1.0, notifier);

    // hold S-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKSlh === 1'b1),
        negedge S &&& (shcheckCKSlh === 1'b1), 1.0, notifier);

    // hold D1-hl CK-lh (!S&!SE)
    $hold(posedge CK &&& (shcheckCKD1lh === 1'b1),
        negedge D1 &&& (shcheckCKD1lh === 1'b1), 1.0, notifier);

    // hold D1-lh CK-lh (!S&!SE)
    $hold(posedge CK &&& (shcheckCKD1lh === 1'b1),
        posedge D1 &&& (shcheckCKD1lh === 1'b1), 1.0, notifier);

    // hold D2-hl CK-lh (S&!SE)
    $hold(posedge CK &&& (shcheckCKD2lh === 1'b1),
        negedge D2 &&& (shcheckCKD2lh === 1'b1), 1.0, notifier);

    // hold D2-lh CK-lh (S&!SE)
    $hold(posedge CK &&& (shcheckCKD2lh === 1'b1),
        posedge D2 &&& (shcheckCKD2lh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HSDFMQM8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:06:24 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HSDFQM1N(D, SD, SE, CK, Q);
  input D, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(shcheckCKDlh, SE);

    buf SMC_I5(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HSDFQM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:06:27 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HSDFQM2N(D, SD, SE, CK, Q);
  input D, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(shcheckCKDlh, SE);

    buf SMC_I5(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HSDFQM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:06:27 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HSDFQM4N(D, SD, SE, CK, Q);
  input D, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(shcheckCKDlh, SE);

    buf SMC_I5(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HSDFQM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:12:41 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HSDFQM8N(D, SD, SE, CK, Q);
  input D, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(shcheckCKDlh, SE);

    buf SMC_I5(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HSDFQM8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:07:56 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HSDFQRM1N(D, RB, SD, SE, CK, Q);
  input D, RB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKDlh, RB, SE_bar);

    and SMC_I6(shcheckCKSDlh, RB, SE);

    buf SMC_I7(shcheckCKSElh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (RB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (RB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (RB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh (RB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (RB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (RB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 1.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HSDFQRM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:10:18 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HSDFQRM2N(D, RB, SD, SE, CK, Q);
  input D, RB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKDlh, RB, SE_bar);

    and SMC_I6(shcheckCKSDlh, RB, SE);

    buf SMC_I7(shcheckCKSElh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (RB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (RB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (RB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh (RB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (RB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (RB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 1.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HSDFQRM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:09:47 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HSDFQRM4N(D, RB, SD, SE, CK, Q);
  input D, RB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKDlh, RB, SE_bar);

    and SMC_I6(shcheckCKSDlh, RB, SE);

    buf SMC_I7(shcheckCKSElh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (RB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (RB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (RB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh (RB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (RB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (RB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 1.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HSDFQRM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:12:31 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HSDFQRM8N(D, RB, SD, SE, CK, Q);
  input D, RB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKDlh, RB, SE_bar);

    and SMC_I6(shcheckCKSDlh, RB, SE);

    buf SMC_I7(shcheckCKSElh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (RB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (RB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (RB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh (RB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (RB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (RB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 1.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HSDFQRM8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:13:30 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HSDFQRSM1N(D, RB, SB, SD, SE, CK, Q);
  input D, RB, SB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(SB));

  `else // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKDlh, RB, SB, SE_bar);

    buf SMC_I6(shcheckCKRBlh, SB);

    buf SMC_I7(shcheckCKSBlh, RB);

    and SMC_I8(shcheckCKSDlh, RB, SB, SE);

    and SMC_I9(shcheckCKSElh, RB, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (RB&SB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (RB&SB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SB-lh RB-lh ()
    $setup(posedge SB, posedge RB, 1.0, notifier);

    // setup SE-hl CK-lh (RB&SB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (RB&SB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (RB&SB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (RB&SB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB&SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB&SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SB-lh RB-lh ()
    $hold(posedge RB, posedge SB, 1.0, notifier);

    // hold SE-hl CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (RB&SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (RB&SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh (SB)
    $recovery(posedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh (RB)
    $recovery(posedge SB &&& (shcheckCKSBlh === 1'b1),
        posedge CK &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // removal RB-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        posedge RB &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // removal SB-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSBlh === 1'b1),
        posedge SB &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HSDFQRSM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:12:10 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HSDFQRSM2N(D, RB, SB, SD, SE, CK, Q);
  input D, RB, SB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(SB));

  `else // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKDlh, RB, SB, SE_bar);

    buf SMC_I6(shcheckCKRBlh, SB);

    buf SMC_I7(shcheckCKSBlh, RB);

    and SMC_I8(shcheckCKSDlh, RB, SB, SE);

    and SMC_I9(shcheckCKSElh, RB, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (RB&SB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (RB&SB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SB-lh RB-lh ()
    $setup(posedge SB, posedge RB, 1.0, notifier);

    // setup SE-hl CK-lh (RB&SB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (RB&SB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (RB&SB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (RB&SB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB&SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB&SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SB-lh RB-lh ()
    $hold(posedge RB, posedge SB, 1.0, notifier);

    // hold SE-hl CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (RB&SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (RB&SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh (SB)
    $recovery(posedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh (RB)
    $recovery(posedge SB &&& (shcheckCKSBlh === 1'b1),
        posedge CK &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // removal RB-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        posedge RB &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // removal SB-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSBlh === 1'b1),
        posedge SB &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HSDFQRSM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:14:54 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HSDFQRSM4N(D, RB, SB, SD, SE, CK, Q);
  input D, RB, SB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(SB));

  `else // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKDlh, RB, SB, SE_bar);

    buf SMC_I6(shcheckCKRBlh, SB);

    buf SMC_I7(shcheckCKSBlh, RB);

    and SMC_I8(shcheckCKSDlh, RB, SB, SE);

    and SMC_I9(shcheckCKSElh, RB, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (RB&SB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (RB&SB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SB-lh RB-lh ()
    $setup(posedge SB, posedge RB, 1.0, notifier);

    // setup SE-hl CK-lh (RB&SB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (RB&SB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (RB&SB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (RB&SB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB&SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB&SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SB-lh RB-lh ()
    $hold(posedge RB, posedge SB, 1.0, notifier);

    // hold SE-hl CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (RB&SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (RB&SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh (SB)
    $recovery(posedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh (RB)
    $recovery(posedge SB &&& (shcheckCKSBlh === 1'b1),
        posedge CK &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // removal RB-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        posedge RB &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // removal SB-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSBlh === 1'b1),
        posedge SB &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HSDFQRSM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:06:38 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HSDFQRSM8N(D, RB, SB, SD, SE, CK, Q);
  input D, RB, SB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(SB));

  `else // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKDlh, RB, SB, SE_bar);

    buf SMC_I6(shcheckCKRBlh, SB);

    buf SMC_I7(shcheckCKSBlh, RB);

    and SMC_I8(shcheckCKSDlh, RB, SB, SE);

    and SMC_I9(shcheckCKSElh, RB, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (RB&SB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (RB&SB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SB-lh RB-lh ()
    $setup(posedge SB, posedge RB, 1.0, notifier);

    // setup SE-hl CK-lh (RB&SB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (RB&SB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (RB&SB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (RB&SB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB&SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB&SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SB-lh RB-lh ()
    $hold(posedge RB, posedge SB, 1.0, notifier);

    // hold SE-hl CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (RB&SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (RB&SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh (SB)
    $recovery(posedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh (RB)
    $recovery(posedge SB &&& (shcheckCKSBlh === 1'b1),
        posedge CK &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // removal RB-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        posedge RB &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // removal SB-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSBlh === 1'b1),
        posedge SB &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HSDFQRSM8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:06:41 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HSDFQSM1N(D, SB, SD, SE, CK, Q);
  input D, SB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(SB));

  `else // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(SB), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKDlh, SB, SE_bar);

    and SMC_I6(shcheckCKSDlh, SB, SE);

    buf SMC_I7(shcheckCKSElh, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (SB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (SB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (SB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh (SB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (SB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 1.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HSDFQSM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:07:51 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HSDFQSM2N(D, SB, SD, SE, CK, Q);
  input D, SB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(SB));

  `else // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(SB), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKDlh, SB, SE_bar);

    and SMC_I6(shcheckCKSDlh, SB, SE);

    buf SMC_I7(shcheckCKSElh, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (SB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (SB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (SB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh (SB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (SB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 1.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HSDFQSM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:12:13 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HSDFQSM4N(D, SB, SD, SE, CK, Q);
  input D, SB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(SB));

  `else // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(SB), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKDlh, SB, SE_bar);

    and SMC_I6(shcheckCKSDlh, SB, SE);

    buf SMC_I7(shcheckCKSElh, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (SB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (SB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (SB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh (SB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (SB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 1.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HSDFQSM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:13:34 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module HSDFQSM8N(D, SB, SD, SE, CK, Q);
  input D, SB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(SB));

  `else // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(SB), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKDlh, SB, SE_bar);

    and SMC_I6(shcheckCKSDlh, SB, SE);

    buf SMC_I7(shcheckCKSElh, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (SB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (SB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (SB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh (SB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (SB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 1.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // HSDFQSM8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:08:45 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module INVM0N(A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // INVM0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:14:02 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module INVM10N(A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // INVM10N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:13:48 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module INVM12N(A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // INVM12N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:08:07 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module INVM14N(A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // INVM14N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:08:06 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module INVM16N(A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // INVM16N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:08:08 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module INVM18N(A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // INVM18N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:08:10 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module INVM1N(A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // INVM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:09:43 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module INVM20N(A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // INVM20N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:10:34 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module INVM2N(A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // INVM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:13:16 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module INVM3N(A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // INVM3N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:07:28 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module INVM4N(A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // INVM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:13:42 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module INVM5N(A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // INVM5N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:12:50 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module INVM6N(A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // INVM6N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:14:01 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module INVM8N(A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // INVM8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:09:56 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LACM0N(D, GB, Q, QB);
  input D, GB;
  output Q, QB;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, GB);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc D --> Q
    (D => Q) = (1.0, 1.0);

    // arc D --> QB
    (D => QB) = (1.0, 1.0);

    // arc GB --> Q
    (negedge GB => ( Q +: D )) = (1.0, 1.0);

    // arc GB --> QB
    (negedge GB => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl GB-lh ()
    $setup(negedge D, posedge GB, 1.0, notifier);

    // setup D-lh GB-lh ()
    $setup(posedge D, posedge GB, 1.0, notifier);

    // hold D-hl GB-lh ()
    $hold(posedge GB, negedge D, 1.0, notifier);

    // hold D-lh GB-lh ()
    $hold(posedge GB, posedge D, 1.0, notifier);

    // mpw GB-lh NS-lh ()
    $width(posedge GB, 1.0, 0, notifier);

    // mpw GB-hl NS-hl ()
    $width(negedge GB, 1.0, 0, notifier);

    $period( posedge GB, 0, notifier );
    $period( negedge GB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LACM0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:14:03 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LACM1N(D, GB, Q, QB);
  input D, GB;
  output Q, QB;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, GB);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc D --> Q
    (D => Q) = (1.0, 1.0);

    // arc D --> QB
    (D => QB) = (1.0, 1.0);

    // arc GB --> Q
    (negedge GB => ( Q +: D )) = (1.0, 1.0);

    // arc GB --> QB
    (negedge GB => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl GB-lh ()
    $setup(negedge D, posedge GB, 1.0, notifier);

    // setup D-lh GB-lh ()
    $setup(posedge D, posedge GB, 1.0, notifier);

    // hold D-hl GB-lh ()
    $hold(posedge GB, negedge D, 1.0, notifier);

    // hold D-lh GB-lh ()
    $hold(posedge GB, posedge D, 1.0, notifier);

    // mpw GB-lh NS-lh ()
    $width(posedge GB, 1.0, 0, notifier);

    // mpw GB-hl NS-hl ()
    $width(negedge GB, 1.0, 0, notifier);

    $period( posedge GB, 0, notifier );
    $period( negedge GB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LACM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:06:56 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LACM2N(D, GB, Q, QB);
  input D, GB;
  output Q, QB;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, GB);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc D --> Q
    (D => Q) = (1.0, 1.0);

    // arc D --> QB
    (D => QB) = (1.0, 1.0);

    // arc GB --> Q
    (negedge GB => ( Q +: D )) = (1.0, 1.0);

    // arc GB --> QB
    (negedge GB => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl GB-lh ()
    $setup(negedge D, posedge GB, 1.0, notifier);

    // setup D-lh GB-lh ()
    $setup(posedge D, posedge GB, 1.0, notifier);

    // hold D-hl GB-lh ()
    $hold(posedge GB, negedge D, 1.0, notifier);

    // hold D-lh GB-lh ()
    $hold(posedge GB, posedge D, 1.0, notifier);

    // mpw GB-lh NS-lh ()
    $width(posedge GB, 1.0, 0, notifier);

    // mpw GB-hl NS-hl ()
    $width(negedge GB, 1.0, 0, notifier);

    $period( posedge GB, 0, notifier );
    $period( negedge GB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LACM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:08:11 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LACM4N(D, GB, Q, QB);
  input D, GB;
  output Q, QB;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, GB);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc D --> Q
    (D => Q) = (1.0, 1.0);

    // arc D --> QB
    (D => QB) = (1.0, 1.0);

    // arc GB --> Q
    (negedge GB => ( Q +: D )) = (1.0, 1.0);

    // arc GB --> QB
    (negedge GB => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl GB-lh ()
    $setup(negedge D, posedge GB, 1.0, notifier);

    // setup D-lh GB-lh ()
    $setup(posedge D, posedge GB, 1.0, notifier);

    // hold D-hl GB-lh ()
    $hold(posedge GB, negedge D, 1.0, notifier);

    // hold D-lh GB-lh ()
    $hold(posedge GB, posedge D, 1.0, notifier);

    // mpw GB-lh NS-lh ()
    $width(posedge GB, 1.0, 0, notifier);

    // mpw GB-hl NS-hl ()
    $width(negedge GB, 1.0, 0, notifier);

    $period( posedge GB, 0, notifier );
    $period( negedge GB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LACM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:12:29 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LACRSM0N(D, RB, SB, GB, Q, QB);
  input D, RB, SB, GB;
  output Q, QB;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, GB);

    inv_clr0 SMC_I1(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ));

  `ifdef functional // functional //
    ldlatch_p1 SMC_I3(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(RB),
        .preset(SB));

  `else // functional //
    ldlatch_p1 SMC_I3(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(RB),
        .preset(SB), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I5(Q, SMC_IQ);

    buf SMC_I6(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I7(shcheckGBDlh, RB, SB);

    buf SMC_I8(shcheckGBRBlh, SB);

    buf SMC_I9(shcheckGBSBlh, RB);

    buf SMC_I10(shcheckRBSBlh, GB);


  specify


    // arc D --> Q
    (D => Q) = (1.0, 1.0);

    // arc D --> QB
    (D => QB) = (1.0, 1.0);

    // arc GB --> Q
    (negedge GB => ( Q +: D )) = (1.0, 1.0);

    // arc GB --> QB
    (negedge GB => ( QB +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl GB-lh (RB&SB)
    $setup(negedge D &&& (shcheckGBDlh === 1'b1),
        posedge GB &&& (shcheckGBDlh === 1'b1), 1.0, notifier);

    // setup D-lh GB-lh (RB&SB)
    $setup(posedge D &&& (shcheckGBDlh === 1'b1),
        posedge GB &&& (shcheckGBDlh === 1'b1), 1.0, notifier);

    // setup SB-lh RB-lh (GB)
    $setup(posedge SB &&& (shcheckRBSBlh === 1'b1),
        posedge RB &&& (shcheckRBSBlh === 1'b1), 1.0, notifier);

    // hold D-hl GB-lh (RB&SB)
    $hold(posedge GB &&& (shcheckGBDlh === 1'b1),
        negedge D &&& (shcheckGBDlh === 1'b1), 1.0, notifier);

    // hold D-lh GB-lh (RB&SB)
    $hold(posedge GB &&& (shcheckGBDlh === 1'b1),
        posedge D &&& (shcheckGBDlh === 1'b1), 1.0, notifier);

    // hold SB-lh RB-lh (GB)
    $hold(posedge RB &&& (shcheckRBSBlh === 1'b1),
        posedge SB &&& (shcheckRBSBlh === 1'b1), 1.0, notifier);

    // recovery RB-lh GB-lh (SB)
    $recovery(posedge RB &&& (shcheckGBRBlh === 1'b1),
        posedge GB &&& (shcheckGBRBlh === 1'b1), 1.0, notifier);

    // recovery SB-lh GB-lh (RB)
    $recovery(posedge SB &&& (shcheckGBSBlh === 1'b1),
        posedge GB &&& (shcheckGBSBlh === 1'b1), 1.0, notifier);

    // removal RB-lh GB-lh (SB)
    $hold(posedge GB &&& (shcheckGBRBlh === 1'b1),
        posedge RB &&& (shcheckGBRBlh === 1'b1), 1.0, notifier);

    // removal SB-lh GB-lh (RB)
    $hold(posedge GB &&& (shcheckGBSBlh === 1'b1),
        posedge SB &&& (shcheckGBSBlh === 1'b1), 1.0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    // mpw GB-hl NS-hl ()
    $width(negedge GB, 1.0, 0, notifier);

    // mpw GB-lh NS-lh ()
    $width(posedge GB, 1.0, 0, notifier);

    $period( posedge GB, 0, notifier );
    $period( negedge GB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LACRSM0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:07:41 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LACRSM1N(D, RB, SB, GB, Q, QB);
  input D, RB, SB, GB;
  output Q, QB;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, GB);

    inv_clr0 SMC_I1(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ));

  `ifdef functional // functional //
    ldlatch_p1 SMC_I3(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(RB),
        .preset(SB));

  `else // functional //
    ldlatch_p1 SMC_I3(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(RB),
        .preset(SB), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I5(Q, SMC_IQ);

    buf SMC_I6(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I7(shcheckGBDlh, RB, SB);

    buf SMC_I8(shcheckGBRBlh, SB);

    buf SMC_I9(shcheckGBSBlh, RB);

    buf SMC_I10(shcheckRBSBlh, GB);


  specify


    // arc D --> Q
    (D => Q) = (1.0, 1.0);

    // arc D --> QB
    (D => QB) = (1.0, 1.0);

    // arc GB --> Q
    (negedge GB => ( Q +: D )) = (1.0, 1.0);

    // arc GB --> QB
    (negedge GB => ( QB +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl GB-lh (RB&SB)
    $setup(negedge D &&& (shcheckGBDlh === 1'b1),
        posedge GB &&& (shcheckGBDlh === 1'b1), 1.0, notifier);

    // setup D-lh GB-lh (RB&SB)
    $setup(posedge D &&& (shcheckGBDlh === 1'b1),
        posedge GB &&& (shcheckGBDlh === 1'b1), 1.0, notifier);

    // setup SB-lh RB-lh (GB)
    $setup(posedge SB &&& (shcheckRBSBlh === 1'b1),
        posedge RB &&& (shcheckRBSBlh === 1'b1), 1.0, notifier);

    // hold D-hl GB-lh (RB&SB)
    $hold(posedge GB &&& (shcheckGBDlh === 1'b1),
        negedge D &&& (shcheckGBDlh === 1'b1), 1.0, notifier);

    // hold D-lh GB-lh (RB&SB)
    $hold(posedge GB &&& (shcheckGBDlh === 1'b1),
        posedge D &&& (shcheckGBDlh === 1'b1), 1.0, notifier);

    // hold SB-lh RB-lh (GB)
    $hold(posedge RB &&& (shcheckRBSBlh === 1'b1),
        posedge SB &&& (shcheckRBSBlh === 1'b1), 1.0, notifier);

    // recovery RB-lh GB-lh (SB)
    $recovery(posedge RB &&& (shcheckGBRBlh === 1'b1),
        posedge GB &&& (shcheckGBRBlh === 1'b1), 1.0, notifier);

    // recovery SB-lh GB-lh (RB)
    $recovery(posedge SB &&& (shcheckGBSBlh === 1'b1),
        posedge GB &&& (shcheckGBSBlh === 1'b1), 1.0, notifier);

    // removal RB-lh GB-lh (SB)
    $hold(posedge GB &&& (shcheckGBRBlh === 1'b1),
        posedge RB &&& (shcheckGBRBlh === 1'b1), 1.0, notifier);

    // removal SB-lh GB-lh (RB)
    $hold(posedge GB &&& (shcheckGBSBlh === 1'b1),
        posedge SB &&& (shcheckGBSBlh === 1'b1), 1.0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    // mpw GB-hl NS-hl ()
    $width(negedge GB, 1.0, 0, notifier);

    // mpw GB-lh NS-lh ()
    $width(posedge GB, 1.0, 0, notifier);

    $period( posedge GB, 0, notifier );
    $period( negedge GB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LACRSM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:14:14 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LACRSM2N(D, RB, SB, GB, Q, QB);
  input D, RB, SB, GB;
  output Q, QB;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, GB);

    inv_clr0 SMC_I1(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ));

  `ifdef functional // functional //
    ldlatch_p1 SMC_I3(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(RB),
        .preset(SB));

  `else // functional //
    ldlatch_p1 SMC_I3(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(RB),
        .preset(SB), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I5(Q, SMC_IQ);

    buf SMC_I6(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I7(shcheckGBDlh, RB, SB);

    buf SMC_I8(shcheckGBRBlh, SB);

    buf SMC_I9(shcheckGBSBlh, RB);

    buf SMC_I10(shcheckRBSBlh, GB);


  specify


    // arc D --> Q
    (D => Q) = (1.0, 1.0);

    // arc D --> QB
    (D => QB) = (1.0, 1.0);

    // arc GB --> Q
    (negedge GB => ( Q +: D )) = (1.0, 1.0);

    // arc GB --> QB
    (negedge GB => ( QB +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl GB-lh (RB&SB)
    $setup(negedge D &&& (shcheckGBDlh === 1'b1),
        posedge GB &&& (shcheckGBDlh === 1'b1), 1.0, notifier);

    // setup D-lh GB-lh (RB&SB)
    $setup(posedge D &&& (shcheckGBDlh === 1'b1),
        posedge GB &&& (shcheckGBDlh === 1'b1), 1.0, notifier);

    // setup SB-lh RB-lh (GB)
    $setup(posedge SB &&& (shcheckRBSBlh === 1'b1),
        posedge RB &&& (shcheckRBSBlh === 1'b1), 1.0, notifier);

    // hold D-hl GB-lh (RB&SB)
    $hold(posedge GB &&& (shcheckGBDlh === 1'b1),
        negedge D &&& (shcheckGBDlh === 1'b1), 1.0, notifier);

    // hold D-lh GB-lh (RB&SB)
    $hold(posedge GB &&& (shcheckGBDlh === 1'b1),
        posedge D &&& (shcheckGBDlh === 1'b1), 1.0, notifier);

    // hold SB-lh RB-lh (GB)
    $hold(posedge RB &&& (shcheckRBSBlh === 1'b1),
        posedge SB &&& (shcheckRBSBlh === 1'b1), 1.0, notifier);

    // recovery RB-lh GB-lh (SB)
    $recovery(posedge RB &&& (shcheckGBRBlh === 1'b1),
        posedge GB &&& (shcheckGBRBlh === 1'b1), 1.0, notifier);

    // recovery SB-lh GB-lh (RB)
    $recovery(posedge SB &&& (shcheckGBSBlh === 1'b1),
        posedge GB &&& (shcheckGBSBlh === 1'b1), 1.0, notifier);

    // removal RB-lh GB-lh (SB)
    $hold(posedge GB &&& (shcheckGBRBlh === 1'b1),
        posedge RB &&& (shcheckGBRBlh === 1'b1), 1.0, notifier);

    // removal SB-lh GB-lh (RB)
    $hold(posedge GB &&& (shcheckGBSBlh === 1'b1),
        posedge SB &&& (shcheckGBSBlh === 1'b1), 1.0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    // mpw GB-hl NS-hl ()
    $width(negedge GB, 1.0, 0, notifier);

    // mpw GB-lh NS-lh ()
    $width(posedge GB, 1.0, 0, notifier);

    $period( posedge GB, 0, notifier );
    $period( negedge GB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LACRSM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:07:53 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LACRSM4N(D, RB, SB, GB, Q, QB);
  input D, RB, SB, GB;
  output Q, QB;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, GB);

    inv_clr0 SMC_I1(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ));

  `ifdef functional // functional //
    ldlatch_p1 SMC_I3(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(RB),
        .preset(SB));

  `else // functional //
    ldlatch_p1 SMC_I3(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(RB),
        .preset(SB), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I5(Q, SMC_IQ);

    buf SMC_I6(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I7(shcheckGBDlh, RB, SB);

    buf SMC_I8(shcheckGBRBlh, SB);

    buf SMC_I9(shcheckGBSBlh, RB);

    buf SMC_I10(shcheckRBSBlh, GB);


  specify


    // arc D --> Q
    (D => Q) = (1.0, 1.0);

    // arc D --> QB
    (D => QB) = (1.0, 1.0);

    // arc GB --> Q
    (negedge GB => ( Q +: D )) = (1.0, 1.0);

    // arc GB --> QB
    (negedge GB => ( QB +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl GB-lh (RB&SB)
    $setup(negedge D &&& (shcheckGBDlh === 1'b1),
        posedge GB &&& (shcheckGBDlh === 1'b1), 1.0, notifier);

    // setup D-lh GB-lh (RB&SB)
    $setup(posedge D &&& (shcheckGBDlh === 1'b1),
        posedge GB &&& (shcheckGBDlh === 1'b1), 1.0, notifier);

    // setup SB-lh RB-lh (GB)
    $setup(posedge SB &&& (shcheckRBSBlh === 1'b1),
        posedge RB &&& (shcheckRBSBlh === 1'b1), 1.0, notifier);

    // hold D-hl GB-lh (RB&SB)
    $hold(posedge GB &&& (shcheckGBDlh === 1'b1),
        negedge D &&& (shcheckGBDlh === 1'b1), 1.0, notifier);

    // hold D-lh GB-lh (RB&SB)
    $hold(posedge GB &&& (shcheckGBDlh === 1'b1),
        posedge D &&& (shcheckGBDlh === 1'b1), 1.0, notifier);

    // hold SB-lh RB-lh (GB)
    $hold(posedge RB &&& (shcheckRBSBlh === 1'b1),
        posedge SB &&& (shcheckRBSBlh === 1'b1), 1.0, notifier);

    // recovery RB-lh GB-lh (SB)
    $recovery(posedge RB &&& (shcheckGBRBlh === 1'b1),
        posedge GB &&& (shcheckGBRBlh === 1'b1), 1.0, notifier);

    // recovery SB-lh GB-lh (RB)
    $recovery(posedge SB &&& (shcheckGBSBlh === 1'b1),
        posedge GB &&& (shcheckGBSBlh === 1'b1), 1.0, notifier);

    // removal RB-lh GB-lh (SB)
    $hold(posedge GB &&& (shcheckGBRBlh === 1'b1),
        posedge RB &&& (shcheckGBRBlh === 1'b1), 1.0, notifier);

    // removal SB-lh GB-lh (RB)
    $hold(posedge GB &&& (shcheckGBSBlh === 1'b1),
        posedge SB &&& (shcheckGBSBlh === 1'b1), 1.0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    // mpw GB-hl NS-hl ()
    $width(negedge GB, 1.0, 0, notifier);

    // mpw GB-lh NS-lh ()
    $width(posedge GB, 1.0, 0, notifier);

    $period( posedge GB, 0, notifier );
    $period( negedge GB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LACRSM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:12:15 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEM12N(E, CK, GCK);
  input E, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I3(GCK, CK, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
  specify


    // arc CK --> GCK
    (CK => GCK) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCEM12N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:10:08 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEM16N(E, CK, GCK);
  input E, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I3(GCK, CK, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
  specify


    // arc CK --> GCK
    (CK => GCK) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCEM16N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:11:48 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEM20N(E, CK, GCK);
  input E, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I3(GCK, CK, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> GCK
    (CK => GCK) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCEM20N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:14:15 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEM2N(E, CK, GCK);
  input E, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I3(GCK, CK, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
  specify


    // arc CK --> GCK
    (CK => GCK) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCEM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:08:13 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEM3N(E, CK, GCK);
  input E, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I3(GCK, CK, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
  specify


    // arc CK --> GCK
    (CK => GCK) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCEM3N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:13:44 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEM4N(E, CK, GCK);
  input E, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I3(GCK, CK, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
  specify


    // arc CK --> GCK
    (CK => GCK) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCEM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:14:15 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEM6N(E, CK, GCK);
  input E, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I3(GCK, CK, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
  specify


    // arc CK --> GCK
    (CK => GCK) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCEM6N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:10:39 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEM8N(E, CK, GCK);
  input E, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I3(GCK, CK, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
  specify


    // arc CK --> GCK
    (CK => GCK) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCEM8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:10:23 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEPM12N(E, SE, CK, GCK);
  input E, SE, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I3(OUT0, CK, SE);
    and SMC_I4(OUT1, CK, SMC_IQ);
    or SMC_I5(GCK, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(shcheckCKSElh, SE);

  specify


    // arc CK --> GCK
    (CK => GCK) = (1.0, 1.0);

    // arc SE --> GCK
    (SE => GCK) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // nochange_setup SE-lh CK-lh (!E)
    $nochange(posedge CK, posedge SE &&& (E===1'b0), 1.0, 1.0);

    // nochange_setup SE-lh CK-lh (E)
    $nochange(posedge CK, posedge SE &&& (E===1'b1), 1.0, 1.0);

    // nochange_setup SE-hl CK-lh (!E)
    $nochange(posedge CK, negedge SE &&& (shcheckCKSElh===1'b1), 1.0, 1.0);

    // nochange_setup SE-hl CK-lh (E)
    $nochange(posedge CK, negedge SE &&& (E===1'b1), 1.0, 1.0);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCEPM12N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:08:08 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEPM16N(E, SE, CK, GCK);
  input E, SE, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I3(OUT0, CK, SE);
    and SMC_I4(OUT1, CK, SMC_IQ);
    or SMC_I5(GCK, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(shcheckCKSElh, SE);

  specify


    // arc CK --> GCK
    (CK => GCK) = (1.0, 1.0);

    // arc SE --> GCK
    (SE => GCK) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // nochange_setup SE-lh CK-lh (!E)
    $nochange(posedge CK, posedge SE &&& (E===1'b0), 1.0, 1.0);

    // nochange_setup SE-lh CK-lh (E)
    $nochange(posedge CK, posedge SE &&& (E===1'b1), 1.0, 1.0);

    // nochange_setup SE-hl CK-lh (!E)
    $nochange(posedge CK, negedge SE &&& (shcheckCKSElh===1'b1), 1.0, 1.0);

    // nochange_setup SE-hl CK-lh (E)
    $nochange(posedge CK, negedge SE &&& (E===1'b1), 1.0, 1.0);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCEPM16N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:14:29 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEPM20N(E, SE, CK, GCK);
  input E, SE, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I3(OUT0, CK, SE);
    and SMC_I4(OUT1, CK, SMC_IQ);
    or SMC_I5(GCK, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(shcheckCKSElh, SE);

  specify


    // arc CK --> GCK
    (CK => GCK) = (1.0, 1.0);

    // arc SE --> GCK
    (SE => GCK) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // nochange_setup SE-lh CK-lh (!E)
    $nochange(posedge CK, posedge SE &&& (E===1'b0), 1.0, 1.0);

    // nochange_setup SE-lh CK-lh (E)
    $nochange(posedge CK, posedge SE &&& (E===1'b1), 1.0, 1.0);

    // nochange_setup SE-hl CK-lh (!E)
    $nochange(posedge CK, negedge SE &&& (shcheckCKSElh===1'b1), 1.0, 1.0);

    // nochange_setup SE-hl CK-lh (E)
    $nochange(posedge CK, negedge SE &&& (E===1'b1), 1.0, 1.0);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCEPM20N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:12:03 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEPM2N(E, SE, CK, GCK);
  input E, SE, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I3(OUT0, CK, SE);
    and SMC_I4(OUT1, CK, SMC_IQ);
    or SMC_I5(GCK, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(shcheckCKSElh, SE);

  specify


    // arc CK --> GCK
    (CK => GCK) = (1.0, 1.0);

    // arc SE --> GCK
    (SE => GCK) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // nochange_setup SE-lh CK-lh (!E)
    $nochange(posedge CK, posedge SE &&& (E===1'b0), 1.0, 1.0);

    // nochange_setup SE-lh CK-lh (E)
    $nochange(posedge CK, posedge SE &&& (E===1'b1), 1.0, 1.0);

    // nochange_setup SE-hl CK-lh (!E)
    $nochange(posedge CK, negedge SE &&& (shcheckCKSElh===1'b1), 1.0, 1.0);

    // nochange_setup SE-hl CK-lh (E)
    $nochange(posedge CK, negedge SE &&& (E===1'b1), 1.0, 1.0);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify
  
  `endif // functional //
endmodule     // LAGCEPM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:12:30 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEPM3N(E, SE, CK, GCK);
  input E, SE, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I3(OUT0, CK, SE);
    and SMC_I4(OUT1, CK, SMC_IQ);
    or SMC_I5(GCK, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(shcheckCKSElh, SE);

  specify


    // arc CK --> GCK
    (CK => GCK) = (1.0, 1.0);

    // arc SE --> GCK
    (SE => GCK) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // nochange_setup SE-lh CK-lh (!E)
    $nochange(posedge CK, posedge SE &&& (E===1'b0), 1.0, 1.0);

    // nochange_setup SE-lh CK-lh (E)
    $nochange(posedge CK, posedge SE &&& (E===1'b1), 1.0, 1.0);

    // nochange_setup SE-hl CK-lh (!E)
    $nochange(posedge CK, negedge SE &&& (shcheckCKSElh===1'b1), 1.0, 1.0);

    // nochange_setup SE-hl CK-lh (E)
    $nochange(posedge CK, negedge SE &&& (E===1'b1), 1.0, 1.0);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCEPM3N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:10:24 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEPM4N(E, SE, CK, GCK);
  input E, SE, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I3(OUT0, CK, SE);
    and SMC_I4(OUT1, CK, SMC_IQ);
    or SMC_I5(GCK, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(shcheckCKSElh, SE);

  specify


    // arc CK --> GCK
    (CK => GCK) = (1.0, 1.0);

    // arc SE --> GCK
    (SE => GCK) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // nochange_setup SE-lh CK-lh (!E)
    $nochange(posedge CK, posedge SE &&& (E===1'b0), 1.0, 1.0);

    // nochange_setup SE-lh CK-lh (E)
    $nochange(posedge CK, posedge SE &&& (E===1'b1), 1.0, 1.0);

    // nochange_setup SE-hl CK-lh (!E)
    $nochange(posedge CK, negedge SE &&& (shcheckCKSElh===1'b1), 1.0, 1.0);

    // nochange_setup SE-hl CK-lh (E)
    $nochange(posedge CK, negedge SE &&& (E===1'b1), 1.0, 1.0);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCEPM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:08:59 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEPM6N(E, SE, CK, GCK);
  input E, SE, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I3(OUT0, CK, SE);
    and SMC_I4(OUT1, CK, SMC_IQ);
    or SMC_I5(GCK, OUT0, OUT1);

  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(shcheckCKSElh, SE);

  specify


    // arc CK --> GCK
    (CK => GCK) = (1.0, 1.0);

    // arc SE --> GCK
    (SE => GCK) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // nochange_setup SE-lh CK-lh (!E)
    $nochange(posedge CK, posedge SE &&& (E===1'b0), 1.0, 1.0);

    // nochange_setup SE-lh CK-lh (E)
    $nochange(posedge CK, posedge SE &&& (E===1'b1), 1.0, 1.0);

    // nochange_setup SE-hl CK-lh (!E)
    $nochange(posedge CK, negedge SE &&& (shcheckCKSElh===1'b1), 1.0, 1.0);

    // nochange_setup SE-hl CK-lh (E)
    $nochange(posedge CK, negedge SE &&& (E===1'b1), 1.0, 1.0);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCEPM6N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:15:20 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEPM8N(E, SE, CK, GCK);
  input E, SE, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I3(OUT0, CK, SE);
    and SMC_I4(OUT1, CK, SMC_IQ);
    or SMC_I5(GCK, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(shcheckCKSElh, SE);

  specify


    // arc CK --> GCK
    (CK => GCK) = (1.0, 1.0);

    // arc SE --> GCK
    (SE => GCK) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // nochange_setup SE-lh CK-lh (!E)
    $nochange(posedge CK, posedge SE &&& (E===1'b0), 1.0, 1.0);

    // nochange_setup SE-lh CK-lh (E)
    $nochange(posedge CK, posedge SE &&& (E===1'b1), 1.0, 1.0);

    // nochange_setup SE-hl CK-lh (!E)
    $nochange(posedge CK, negedge SE &&& (shcheckCKSElh===1'b1), 1.0, 1.0);

    // nochange_setup SE-hl CK-lh (E)
    $nochange(posedge CK, negedge SE &&& (E===1'b1), 1.0, 1.0);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCEPM8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:08:17 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEPOM12N(E, SE, CK, GCK, OBS);
  input E, SE, CK;
  output GCK, OBS;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(OBS, SMC_IQ);

    and SMC_I4(OUT0, CK, SE);
    and SMC_I5(OUT1, CK, SMC_IQ);
    or SMC_I6(GCK, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //


  specify


    // arc CK --> GCK
    (CK => GCK) = (1.0, 1.0);

    // arc CK --> OBS
    ( negedge CK => ( OBS +: CK ) ) = (1.0, 1.0);

    // arc E --> OBS
    (E => OBS) = (1.0, 1.0);

    // arc SE --> GCK
    (SE => GCK) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // nochange_setup E-lh CK-hl ()
    $nochange(negedge CK, posedge E, 1.0, 1.0);

    // nochange_setup E-hl CK-hl ()
    $nochange(negedge CK, negedge E, 1.0, 1.0);

    // nochange_setup SE-lh CK-lh (!E)
    $nochange(posedge CK, posedge SE &&& (E===1'b0), 1.0, 1.0);

    // nochange_setup SE-lh CK-lh (E)
    $nochange(posedge CK, posedge SE &&& (E===1'b1), 1.0, 1.0);

    // nochange_setup SE-hl CK-lh (!E)
    $nochange(posedge CK, negedge SE &&& (E===1'b0), 1.0, 1.0);

    // nochange_setup SE-hl CK-lh (E)
    $nochange(posedge CK, negedge SE &&& (E===1'b1), 1.0, 1.0);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCEPOM12N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:13:49 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEPOM16N(E, SE, CK, GCK, OBS);
  input E, SE, CK;
  output GCK, OBS;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(OBS, SMC_IQ);

    and SMC_I4(OUT0, CK, SE);
    and SMC_I5(OUT1, CK, SMC_IQ);
    or SMC_I6(GCK, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //


  specify


    // arc CK --> GCK
    (CK => GCK) = (1.0, 1.0);

    // arc CK --> OBS
    ( negedge CK => ( OBS +: CK ) ) = (1.0, 1.0);

    // arc E --> OBS
    (E => OBS) = (1.0, 1.0);

    // arc SE --> GCK
    (SE => GCK) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // nochange_setup E-lh CK-hl ()
    $nochange(negedge CK, posedge E, 1.0, 1.0);

    // nochange_setup E-hl CK-hl ()
    $nochange(negedge CK, negedge E, 1.0, 1.0);

    // nochange_setup SE-lh CK-lh (!E)
    $nochange(posedge CK, posedge SE &&& (E===1'b0), 1.0, 1.0);

    // nochange_setup SE-lh CK-lh (E)
    $nochange(posedge CK, posedge SE &&& (E===1'b1), 1.0, 1.0);

    // nochange_setup SE-hl CK-lh (!E)
    $nochange(posedge CK, negedge SE &&& (E===1'b0), 1.0, 1.0);

    // nochange_setup SE-hl CK-lh (E)
    $nochange(posedge CK, negedge SE &&& (E===1'b1), 1.0, 1.0);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCEPOM16N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:14:18 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEPOM20N(E, SE, CK, GCK, OBS);
  input E, SE, CK;
  output GCK, OBS;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(OBS, SMC_IQ);

    and SMC_I4(OUT0, CK, SE);
    and SMC_I5(OUT1, CK, SMC_IQ);
    or SMC_I6(GCK, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //


  specify


    // arc CK --> GCK
    (CK => GCK) = (1.0, 1.0);

    // arc CK --> OBS
    ( negedge CK => ( OBS +: CK ) ) = (1.0, 1.0);

    // arc E --> OBS
    (E => OBS) = (1.0, 1.0);

    // arc SE --> GCK
    (SE => GCK) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // nochange_setup E-lh CK-hl ()
    $nochange(negedge CK, posedge E, 1.0, 1.0);

    // nochange_setup E-hl CK-hl ()
    $nochange(negedge CK, negedge E, 1.0, 1.0);

    // nochange_setup SE-lh CK-lh (!E)
    $nochange(posedge CK, posedge SE &&& (E===1'b0), 1.0, 1.0);

    // nochange_setup SE-lh CK-lh (E)
    $nochange(posedge CK, posedge SE &&& (E===1'b1), 1.0, 1.0);

    // nochange_setup SE-hl CK-lh (!E)
    $nochange(posedge CK, negedge SE &&& (E===1'b0), 1.0, 1.0);

    // nochange_setup SE-hl CK-lh (E)
    $nochange(posedge CK, negedge SE &&& (E===1'b1), 1.0, 1.0);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCEPOM20N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:12:58 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEPOM2N(E, SE, CK, GCK, OBS);
  input E, SE, CK;
  output GCK, OBS;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(OBS, SMC_IQ);

    and SMC_I4(OUT0, CK, SE);
    and SMC_I5(OUT1, CK, SMC_IQ);
    or SMC_I6(GCK, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //


  specify


    // arc CK --> GCK
    (CK => GCK) = (1.0, 1.0);

    // arc CK --> OBS
    ( negedge CK => ( OBS +: CK ) ) = (1.0, 1.0);

    // arc E --> OBS
    (E => OBS) = (1.0, 1.0);

    // arc SE --> GCK
    (SE => GCK) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // nochange_setup E-lh CK-hl ()
    $nochange(negedge CK, posedge E, 1.0, 1.0);

    // nochange_setup E-hl CK-hl ()
    $nochange(negedge CK, negedge E, 1.0, 1.0);

    // nochange_setup SE-lh CK-lh (!E)
    $nochange(posedge CK, posedge SE &&& (E===1'b0), 1.0, 1.0);

    // nochange_setup SE-lh CK-lh (E)
    $nochange(posedge CK, posedge SE &&& (E===1'b1), 1.0, 1.0);

    // nochange_setup SE-hl CK-lh (!E)
    $nochange(posedge CK, negedge SE &&& (E===1'b0), 1.0, 1.0);

    // nochange_setup SE-hl CK-lh (E)
    $nochange(posedge CK, negedge SE &&& (E===1'b1), 1.0, 1.0);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCEPOM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:10:47 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEPOM3N(E, SE, CK, GCK, OBS);
  input E, SE, CK;
  output GCK, OBS;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(OBS, SMC_IQ);

    and SMC_I4(OUT0, CK, SE);
    and SMC_I5(OUT1, CK, SMC_IQ);
    or SMC_I6(GCK, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //


  specify


    // arc CK --> GCK
    (CK => GCK) = (1.0, 1.0);

    // arc CK --> OBS
    ( negedge CK => ( OBS +: CK ) ) = (1.0, 1.0);

    // arc E --> OBS
    (E => OBS) = (1.0, 1.0);

    // arc SE --> GCK
    (SE => GCK) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // nochange_setup E-lh CK-hl ()
    $nochange(negedge CK, posedge E, 1.0, 1.0);

    // nochange_setup E-hl CK-hl ()
    $nochange(negedge CK, negedge E, 1.0, 1.0);

    // nochange_setup SE-lh CK-lh (!E)
    $nochange(posedge CK, posedge SE &&& (E===1'b0), 1.0, 1.0);

    // nochange_setup SE-lh CK-lh (E)
    $nochange(posedge CK, posedge SE &&& (E===1'b1), 1.0, 1.0);

    // nochange_setup SE-hl CK-lh (!E)
    $nochange(posedge CK, negedge SE &&& (E===1'b0), 1.0, 1.0);

    // nochange_setup SE-hl CK-lh (E)
    $nochange(posedge CK, negedge SE &&& (E===1'b1), 1.0, 1.0);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify
  
  `endif // functional //
endmodule     // LAGCEPOM3N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:13:29 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEPOM4N(E, SE, CK, GCK, OBS);
  input E, SE, CK;
  output GCK, OBS;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(OBS, SMC_IQ);

    and SMC_I4(OUT0, CK, SE);
    and SMC_I5(OUT1, CK, SMC_IQ);
    or SMC_I6(GCK, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //


  specify


    // arc CK --> GCK
    (CK => GCK) = (1.0, 1.0);

    // arc CK --> OBS
    ( negedge CK => ( OBS +: CK ) ) = (1.0, 1.0);

    // arc E --> OBS
    (E => OBS) = (1.0, 1.0);

    // arc SE --> GCK
    (SE => GCK) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // nochange_setup E-lh CK-hl ()
    $nochange(negedge CK, posedge E, 1.0, 1.0);

    // nochange_setup E-hl CK-hl ()
    $nochange(negedge CK, negedge E, 1.0, 1.0);

    // nochange_setup SE-lh CK-lh (!E)
    $nochange(posedge CK, posedge SE &&& (E===1'b0), 1.0, 1.0);

    // nochange_setup SE-lh CK-lh (E)
    $nochange(posedge CK, posedge SE &&& (E===1'b1), 1.0, 1.0);

    // nochange_setup SE-hl CK-lh (!E)
    $nochange(posedge CK, negedge SE &&& (E===1'b0), 1.0, 1.0);

    // nochange_setup SE-hl CK-lh (E)
    $nochange(posedge CK, negedge SE &&& (E===1'b1), 1.0, 1.0);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCEPOM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:11:24 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEPOM6N(E, SE, CK, GCK, OBS);
  input E, SE, CK;
  output GCK, OBS;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(OBS, SMC_IQ);

    and SMC_I4(OUT0, CK, SE);
    and SMC_I5(OUT1, CK, SMC_IQ);
    or SMC_I6(GCK, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //


  specify


    // arc CK --> GCK
    (CK => GCK) = (1.0, 1.0);

    // arc CK --> OBS
    ( negedge CK => ( OBS +: CK ) ) = (1.0, 1.0);

    // arc E --> OBS
    (E => OBS) = (1.0, 1.0);

    // arc SE --> GCK
    (SE => GCK) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // nochange_setup E-lh CK-hl ()
    $nochange(negedge CK, posedge E, 1.0, 1.0);

    // nochange_setup E-hl CK-hl ()
    $nochange(negedge CK, negedge E, 1.0, 1.0);

    // nochange_setup SE-lh CK-lh (!E)
    $nochange(posedge CK, posedge SE &&& (E===1'b0), 1.0, 1.0);

    // nochange_setup SE-lh CK-lh (E)
    $nochange(posedge CK, posedge SE &&& (E===1'b1), 1.0, 1.0);

    // nochange_setup SE-hl CK-lh (!E)
    $nochange(posedge CK, negedge SE &&& (E===1'b0), 1.0, 1.0);

    // nochange_setup SE-hl CK-lh (E)
    $nochange(posedge CK, negedge SE &&& (E===1'b1), 1.0, 1.0);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCEPOM6N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:10:39 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEPOM8N(E, SE, CK, GCK, OBS);
  input E, SE, CK;
  output GCK, OBS;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1), 
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(OBS, SMC_IQ);

    and SMC_I4(OUT0, CK, SE);
    and SMC_I5(OUT1, CK, SMC_IQ);
    or SMC_I6(GCK, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //


  specify


    // arc CK --> GCK
    (CK => GCK) = (1.0, 1.0);

    // arc CK --> OBS
    ( negedge CK => ( OBS +: CK ) ) = (1.0, 1.0);

    // arc E --> OBS
    (E => OBS) = (1.0, 1.0);

    // arc SE --> GCK
    (SE => GCK) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // nochange_setup E-lh CK-hl ()
    $nochange(negedge CK, posedge E, 1.0, 1.0);

    // nochange_setup E-hl CK-hl ()
    $nochange(negedge CK, negedge E, 1.0, 1.0);

    // nochange_setup SE-lh CK-lh (!E)
    $nochange(posedge CK, posedge SE &&& (E===1'b0), 1.0, 1.0);

    // nochange_setup SE-lh CK-lh (E)
    $nochange(posedge CK, posedge SE &&& (E===1'b1), 1.0, 1.0);

    // nochange_setup SE-hl CK-lh (!E)
    $nochange(posedge CK, negedge SE &&& (E===1'b0), 1.0, 1.0);

    // nochange_setup SE-hl CK-lh (E)
    $nochange(posedge CK, negedge SE &&& (E===1'b1), 1.0, 1.0);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCEPOM8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:12:46 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCESM12N(E, SE, CK, GCK);
  input E, SE, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

  wire SMC_LD_IN;
    buf SMC_I1(OUT0, E);
    buf SMC_I2(OUT1, SE);
    or SMC_I3(SMC_LD_IN, OUT0, OUT1);

    not SMC_I4(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN), 
          .clear(1'b1), .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN), 
          .clear(1'b1), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I6(GCK, CK, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> GCK
    (CK => GCK) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCESM12N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:08:24 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCESM16N(E, SE, CK, GCK);
  input E, SE, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

  wire SMC_LD_IN;
    buf SMC_I1(OUT0, E);
    buf SMC_I2(OUT1, SE);
    or SMC_I3(SMC_LD_IN, OUT0, OUT1);

    not SMC_I4(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN), 
          .clear(1'b1), .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN), 
          .clear(1'b1), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I6(GCK, CK, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> GCK
    (CK => GCK) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCESM16N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:10:40 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCESM20N(E, SE, CK, GCK);
  input E, SE, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

  wire SMC_LD_IN;
    buf SMC_I1(OUT0, E);
    buf SMC_I2(OUT1, SE);
    or SMC_I3(SMC_LD_IN, OUT0, OUT1);

    not SMC_I4(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN), 
          .clear(1'b1), .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN), 
          .clear(1'b1), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I6(GCK, CK, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> GCK
    (CK => GCK) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCESM20N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:14:45 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCESM2N(E, SE, CK, GCK);
  input E, SE, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

  wire SMC_LD_IN;
    buf SMC_I1(OUT0, E);
    buf SMC_I2(OUT1, SE);
    or SMC_I3(SMC_LD_IN, OUT0, OUT1);

    not SMC_I4(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN), 
          .clear(1'b1), .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN), 
          .clear(1'b1), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I6(GCK, CK, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> GCK
    (CK => GCK) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCESM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:12:19 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCESM3N(E, SE, CK, GCK);
  input E, SE, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

  wire SMC_LD_IN;
    buf SMC_I1(OUT0, E);
    buf SMC_I2(OUT1, SE);
    or SMC_I3(SMC_LD_IN, OUT0, OUT1);

    not SMC_I4(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN), 
          .clear(1'b1), .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN), 
          .clear(1'b1), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I6(GCK, CK, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> GCK
    (CK => GCK) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCESM3N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:10:50 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCESM4N(E, SE, CK, GCK);
  input E, SE, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

  wire SMC_LD_IN;
    buf SMC_I1(OUT0, E);
    buf SMC_I2(OUT1, SE);
    or SMC_I3(SMC_LD_IN, OUT0, OUT1);

    not SMC_I4(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN), 
          .clear(1'b1), .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN), 
          .clear(1'b1), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I6(GCK, CK, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> GCK
    (CK => GCK) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCESM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:13:33 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCESM6N(E, SE, CK, GCK);
  input E, SE, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

  wire SMC_LD_IN;
    buf SMC_I1(OUT0, E);
    buf SMC_I2(OUT1, SE);
    or SMC_I3(SMC_LD_IN, OUT0, OUT1);

    not SMC_I4(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN), 
          .clear(1'b1), .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN), 
          .clear(1'b1), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I6(GCK, CK, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> GCK
    (CK => GCK) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCESM6N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:11:28 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCESM8N(E, SE, CK, GCK);
  input E, SE, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

  wire SMC_LD_IN;
    buf SMC_I1(OUT0, E);
    buf SMC_I2(OUT1, SE);
    or SMC_I3(SMC_LD_IN, OUT0, OUT1);

    not SMC_I4(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN), 
          .clear(1'b1), .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN), 
          .clear(1'b1), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I6(GCK, CK, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> GCK
    (CK => GCK) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCESM8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:09:12 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCESOM12N(E, SE, CK, GCK, OBS);
  input E, SE, CK;
  output GCK, OBS;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

  wire SMC_LD_IN;
    buf SMC_I1(OUT0, E);
    buf SMC_I2(OUT1, SE);
    or SMC_I3(SMC_LD_IN, OUT0, OUT1);

    not SMC_I4(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN), 
          .clear(1'b1), .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN), 
          .clear(1'b1), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I6(GCK, CK, SMC_IQ);

    buf SMC_I7(OBS, E);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> GCK
    (CK => GCK) = (1.0, 1.0);

    // arc E --> OBS
    (E => OBS) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCESOM12N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:10:56 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCESOM16N(E, SE, CK, GCK, OBS);
  input E, SE, CK;
  output GCK, OBS;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

  wire SMC_LD_IN;
    buf SMC_I1(OUT0, E);
    buf SMC_I2(OUT1, SE);
    or SMC_I3(SMC_LD_IN, OUT0, OUT1);

    not SMC_I4(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN), 
          .clear(1'b1), .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN), 
          .clear(1'b1), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I6(GCK, CK, SMC_IQ);

    buf SMC_I7(OBS, E);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> GCK
    (CK => GCK) = (1.0, 1.0);

    // arc E --> OBS
    (E => OBS) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCESOM16N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:15:01 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCESOM20N(E, SE, CK, GCK, OBS);
  input E, SE, CK;
  output GCK, OBS;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

  wire SMC_LD_IN;
    buf SMC_I1(OUT0, E);
    buf SMC_I2(OUT1, SE);
    or SMC_I3(SMC_LD_IN, OUT0, OUT1);

    not SMC_I4(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN), 
          .clear(1'b1), .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN), 
          .clear(1'b1), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I6(GCK, CK, SMC_IQ);

    buf SMC_I7(OBS, E);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> GCK
    (CK => GCK) = (1.0, 1.0);

    // arc E --> OBS
    (E => OBS) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCESOM20N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:15:15 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCESOM2N(E, SE, CK, GCK, OBS);
  input E, SE, CK;
  output GCK, OBS;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

  wire SMC_LD_IN;
    buf SMC_I1(OUT0, E);
    buf SMC_I2(OUT1, SE);
    or SMC_I3(SMC_LD_IN, OUT0, OUT1);

    not SMC_I4(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN), 
          .clear(1'b1), .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN), 
          .clear(1'b1), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I6(GCK, CK, SMC_IQ);

    buf SMC_I7(OBS, E);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> GCK
    (CK => GCK) = (1.0, 1.0);

    // arc E --> OBS
    (E => OBS) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCESOM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:11:09 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCESOM3N(E, SE, CK, GCK, OBS);
  input E, SE, CK;
  output GCK, OBS;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

  wire SMC_LD_IN;
    buf SMC_I1(OUT0, E);
    buf SMC_I2(OUT1, SE);
    or SMC_I3(SMC_LD_IN, OUT0, OUT1);

    not SMC_I4(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN), 
          .clear(1'b1), .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN), 
          .clear(1'b1), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I6(GCK, CK, SMC_IQ);

    buf SMC_I7(OBS, E);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> GCK
    (CK => GCK) = (1.0, 1.0);

    // arc E --> OBS
    (E => OBS) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCESOM3N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:12:49 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCESOM4N(E, SE, CK, GCK, OBS);
  input E, SE, CK;
  output GCK, OBS;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

  wire SMC_LD_IN;
    buf SMC_I1(OUT0, E);
    buf SMC_I2(OUT1, SE);
    or SMC_I3(SMC_LD_IN, OUT0, OUT1);

    not SMC_I4(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN), 
          .clear(1'b1), .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN), 
          .clear(1'b1), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I6(GCK, CK, SMC_IQ);

    buf SMC_I7(OBS, E);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> GCK
    (CK => GCK) = (1.0, 1.0);

    // arc E --> OBS
    (E => OBS) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCESOM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:14:11 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCESOM6N(E, SE, CK, GCK, OBS);
  input E, SE, CK;
  output GCK, OBS;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

  wire SMC_LD_IN;
    buf SMC_I1(OUT0, E);
    buf SMC_I2(OUT1, SE);
    or SMC_I3(SMC_LD_IN, OUT0, OUT1);

    not SMC_I4(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN), 
          .clear(1'b1), .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN), 
          .clear(1'b1), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I6(GCK, CK, SMC_IQ);

    buf SMC_I7(OBS, E);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> GCK
    (CK => GCK) = (1.0, 1.0);

    // arc E --> OBS
    (E => OBS) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCESOM6N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:08:54 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCESOM8N(E, SE, CK, GCK, OBS);
  input E, SE, CK;
  output GCK, OBS;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

  wire SMC_LD_IN;
    buf SMC_I1(OUT0, E);
    buf SMC_I2(OUT1, SE);
    or SMC_I3(SMC_LD_IN, OUT0, OUT1);

    not SMC_I4(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN), 
          .clear(1'b1), .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN), 
          .clear(1'b1), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I6(GCK, CK, SMC_IQ);

    buf SMC_I7(OBS, E);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> GCK
    (CK => GCK) = (1.0, 1.0);

    // arc E --> OBS
    (E => OBS) = (1.0, 1.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 1.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 1.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCESOM8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:08:10 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAM0N(D, G, Q, QB);
  input D, G;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc D --> Q
    (D => Q) = (1.0, 1.0);

    // arc D --> QB
    (D => QB) = (1.0, 1.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (1.0, 1.0);

    // arc G --> QB
    (posedge G => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl G-hl ()
    $setup(negedge D, negedge G, 1.0, notifier);

    // setup D-lh G-hl ()
    $setup(posedge D, negedge G, 1.0, notifier);

    // hold D-hl G-hl ()
    $hold(negedge G, negedge D, 1.0, notifier);

    // hold D-lh G-hl ()
    $hold(negedge G, posedge D, 1.0, notifier);

    // mpw G-hl NS-hl ()
    $width(negedge G, 1.0, 0, notifier);

    // mpw G-lh NS-lh ()
    $width(posedge G, 1.0, 0, notifier);

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAM0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:15:36 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAM1N(D, G, Q, QB);
  input D, G;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc D --> Q
    (D => Q) = (1.0, 1.0);

    // arc D --> QB
    (D => QB) = (1.0, 1.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (1.0, 1.0);

    // arc G --> QB
    (posedge G => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl G-hl ()
    $setup(negedge D, negedge G, 1.0, notifier);

    // setup D-lh G-hl ()
    $setup(posedge D, negedge G, 1.0, notifier);

    // hold D-hl G-hl ()
    $hold(negedge G, negedge D, 1.0, notifier);

    // hold D-lh G-hl ()
    $hold(negedge G, posedge D, 1.0, notifier);

    // mpw G-hl NS-hl ()
    $width(negedge G, 1.0, 0, notifier);

    // mpw G-lh NS-lh ()
    $width(posedge G, 1.0, 0, notifier);

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:13:35 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAM2N(D, G, Q, QB);
  input D, G;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc D --> Q
    (D => Q) = (1.0, 1.0);

    // arc D --> QB
    (D => QB) = (1.0, 1.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (1.0, 1.0);

    // arc G --> QB
    (posedge G => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl G-hl ()
    $setup(negedge D, negedge G, 1.0, notifier);

    // setup D-lh G-hl ()
    $setup(posedge D, negedge G, 1.0, notifier);

    // hold D-hl G-hl ()
    $hold(negedge G, negedge D, 1.0, notifier);

    // hold D-lh G-hl ()
    $hold(negedge G, posedge D, 1.0, notifier);

    // mpw G-hl NS-hl ()
    $width(negedge G, 1.0, 0, notifier);

    // mpw G-lh NS-lh ()
    $width(posedge G, 1.0, 0, notifier);

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:11:31 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAM4N(D, G, Q, QB);
  input D, G;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc D --> Q
    (D => Q) = (1.0, 1.0);

    // arc D --> QB
    (D => QB) = (1.0, 1.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (1.0, 1.0);

    // arc G --> QB
    (posedge G => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl G-hl ()
    $setup(negedge D, negedge G, 1.0, notifier);

    // setup D-lh G-hl ()
    $setup(posedge D, negedge G, 1.0, notifier);

    // hold D-hl G-hl ()
    $hold(negedge G, negedge D, 1.0, notifier);

    // hold D-lh G-hl ()
    $hold(negedge G, posedge D, 1.0, notifier);

    // mpw G-hl NS-hl ()
    $width(negedge G, 1.0, 0, notifier);

    // mpw G-lh NS-lh ()
    $width(posedge G, 1.0, 0, notifier);

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:13:10 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LARSM0N(D, RB, SB, G, Q, QB);
  input D, RB, SB, G;
  output Q, QB;
  reg notifier;

    inv_clr0 SMC_I0(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ));

  `ifdef functional // functional //
    ldlatch_p1 SMC_I2(.q(SMC_IQ), .d(D), .en(G), .clear(RB), .preset(SB));

  `else // functional //
    ldlatch_p1 SMC_I2(.q(SMC_IQ), .d(D), .en(G), .clear(RB), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I6(shcheckGDhl, RB, SB);

    buf SMC_I7(shcheckGRBhl, SB);

    buf SMC_I8(shcheckGSBhl, RB);

    not SMC_I9(shcheckRBSBlh, G);


  specify


    // arc D --> Q
    (D => Q) = (1.0, 1.0);

    // arc D --> QB
    (D => QB) = (1.0, 1.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (1.0, 1.0);

    // arc G --> QB
    (posedge G => ( QB +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl G-hl (RB&SB)
    $setup(negedge D &&& (shcheckGDhl === 1'b1),
        negedge G &&& (shcheckGDhl === 1'b1), 1.0, notifier);

    // setup D-lh G-hl (RB&SB)
    $setup(posedge D &&& (shcheckGDhl === 1'b1),
        negedge G &&& (shcheckGDhl === 1'b1), 1.0, notifier);

    // setup SB-lh RB-lh (!G)
    $setup(posedge SB &&& (shcheckRBSBlh === 1'b1),
        posedge RB &&& (shcheckRBSBlh === 1'b1), 1.0, notifier);

    // hold D-hl G-hl (RB&SB)
    $hold(negedge G &&& (shcheckGDhl === 1'b1),
        negedge D &&& (shcheckGDhl === 1'b1), 1.0, notifier);

    // hold D-lh G-hl (RB&SB)
    $hold(negedge G &&& (shcheckGDhl === 1'b1),
        posedge D &&& (shcheckGDhl === 1'b1), 1.0, notifier);

    // hold SB-lh RB-lh (!G)
    $hold(posedge RB &&& (shcheckRBSBlh === 1'b1),
        posedge SB &&& (shcheckRBSBlh === 1'b1), 1.0, notifier);

    // recovery SB-lh G-hl (RB)
    $recovery(posedge SB &&& (shcheckGSBhl === 1'b1),
        negedge G &&& (shcheckGSBhl === 1'b1), 1.0, notifier);

    // recovery RB-lh G-hl (SB)
    $recovery(posedge RB &&& (shcheckGRBhl === 1'b1),
        negedge G &&& (shcheckGRBhl === 1'b1), 1.0, notifier);

    // removal SB-lh G-hl (RB)
    $hold(negedge G &&& (shcheckGSBhl === 1'b1),
        posedge SB &&& (shcheckGSBhl === 1'b1), 1.0, notifier);

    // removal RB-lh G-hl (SB)
    $hold(negedge G &&& (shcheckGRBhl === 1'b1),
        posedge RB &&& (shcheckGRBhl === 1'b1), 1.0, notifier);

    // mpw G-lh NS-lh ()
    $width(posedge G, 1.0, 0, notifier);

    // mpw G-hl NS-hl ()
    $width(negedge G, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LARSM0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:13:56 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LARSM1N(D, RB, SB, G, Q, QB);
  input D, RB, SB, G;
  output Q, QB;
  reg notifier;

    inv_clr0 SMC_I0(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ));

  `ifdef functional // functional //
    ldlatch_p1 SMC_I2(.q(SMC_IQ), .d(D), .en(G), .clear(RB), .preset(SB));

  `else // functional //
    ldlatch_p1 SMC_I2(.q(SMC_IQ), .d(D), .en(G), .clear(RB), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I6(shcheckGDhl, RB, SB);

    buf SMC_I7(shcheckGRBhl, SB);

    buf SMC_I8(shcheckGSBhl, RB);

    not SMC_I9(shcheckRBSBlh, G);


  specify


    // arc D --> Q
    (D => Q) = (1.0, 1.0);

    // arc D --> QB
    (D => QB) = (1.0, 1.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (1.0, 1.0);

    // arc G --> QB
    (posedge G => ( QB +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl G-hl (RB&SB)
    $setup(negedge D &&& (shcheckGDhl === 1'b1),
        negedge G &&& (shcheckGDhl === 1'b1), 1.0, notifier);

    // setup D-lh G-hl (RB&SB)
    $setup(posedge D &&& (shcheckGDhl === 1'b1),
        negedge G &&& (shcheckGDhl === 1'b1), 1.0, notifier);

    // setup SB-lh RB-lh (!G)
    $setup(posedge SB &&& (shcheckRBSBlh === 1'b1),
        posedge RB &&& (shcheckRBSBlh === 1'b1), 1.0, notifier);

    // hold D-hl G-hl (RB&SB)
    $hold(negedge G &&& (shcheckGDhl === 1'b1),
        negedge D &&& (shcheckGDhl === 1'b1), 1.0, notifier);

    // hold D-lh G-hl (RB&SB)
    $hold(negedge G &&& (shcheckGDhl === 1'b1),
        posedge D &&& (shcheckGDhl === 1'b1), 1.0, notifier);

    // hold SB-lh RB-lh (!G)
    $hold(posedge RB &&& (shcheckRBSBlh === 1'b1),
        posedge SB &&& (shcheckRBSBlh === 1'b1), 1.0, notifier);

    // recovery SB-lh G-hl (RB)
    $recovery(posedge SB &&& (shcheckGSBhl === 1'b1),
        negedge G &&& (shcheckGSBhl === 1'b1), 1.0, notifier);

    // recovery RB-lh G-hl (SB)
    $recovery(posedge RB &&& (shcheckGRBhl === 1'b1),
        negedge G &&& (shcheckGRBhl === 1'b1), 1.0, notifier);

    // removal SB-lh G-hl (RB)
    $hold(negedge G &&& (shcheckGSBhl === 1'b1),
        posedge SB &&& (shcheckGSBhl === 1'b1), 1.0, notifier);

    // removal RB-lh G-hl (SB)
    $hold(negedge G &&& (shcheckGRBhl === 1'b1),
        posedge RB &&& (shcheckGRBhl === 1'b1), 1.0, notifier);

    // mpw G-lh NS-lh ()
    $width(posedge G, 1.0, 0, notifier);

    // mpw G-hl NS-hl ()
    $width(negedge G, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LARSM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:14:26 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LARSM2N(D, RB, SB, G, Q, QB);
  input D, RB, SB, G;
  output Q, QB;
  reg notifier;

    inv_clr0 SMC_I0(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ));

  `ifdef functional // functional //
    ldlatch_p1 SMC_I2(.q(SMC_IQ), .d(D), .en(G), .clear(RB), .preset(SB));

  `else // functional //
    ldlatch_p1 SMC_I2(.q(SMC_IQ), .d(D), .en(G), .clear(RB), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I6(shcheckGDhl, RB, SB);

    buf SMC_I7(shcheckGRBhl, SB);

    buf SMC_I8(shcheckGSBhl, RB);

    not SMC_I9(shcheckRBSBlh, G);


  specify


    // arc D --> Q
    (D => Q) = (1.0, 1.0);

    // arc D --> QB
    (D => QB) = (1.0, 1.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (1.0, 1.0);

    // arc G --> QB
    (posedge G => ( QB +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl G-hl (RB&SB)
    $setup(negedge D &&& (shcheckGDhl === 1'b1),
        negedge G &&& (shcheckGDhl === 1'b1), 1.0, notifier);

    // setup D-lh G-hl (RB&SB)
    $setup(posedge D &&& (shcheckGDhl === 1'b1),
        negedge G &&& (shcheckGDhl === 1'b1), 1.0, notifier);

    // setup SB-lh RB-lh (!G)
    $setup(posedge SB &&& (shcheckRBSBlh === 1'b1),
        posedge RB &&& (shcheckRBSBlh === 1'b1), 1.0, notifier);

    // hold D-hl G-hl (RB&SB)
    $hold(negedge G &&& (shcheckGDhl === 1'b1),
        negedge D &&& (shcheckGDhl === 1'b1), 1.0, notifier);

    // hold D-lh G-hl (RB&SB)
    $hold(negedge G &&& (shcheckGDhl === 1'b1),
        posedge D &&& (shcheckGDhl === 1'b1), 1.0, notifier);

    // hold SB-lh RB-lh (!G)
    $hold(posedge RB &&& (shcheckRBSBlh === 1'b1),
        posedge SB &&& (shcheckRBSBlh === 1'b1), 1.0, notifier);

    // recovery SB-lh G-hl (RB)
    $recovery(posedge SB &&& (shcheckGSBhl === 1'b1),
        negedge G &&& (shcheckGSBhl === 1'b1), 1.0, notifier);

    // recovery RB-lh G-hl (SB)
    $recovery(posedge RB &&& (shcheckGRBhl === 1'b1),
        negedge G &&& (shcheckGRBhl === 1'b1), 1.0, notifier);

    // removal SB-lh G-hl (RB)
    $hold(negedge G &&& (shcheckGSBhl === 1'b1),
        posedge SB &&& (shcheckGSBhl === 1'b1), 1.0, notifier);

    // removal RB-lh G-hl (SB)
    $hold(negedge G &&& (shcheckGRBhl === 1'b1),
        posedge RB &&& (shcheckGRBhl === 1'b1), 1.0, notifier);

    // mpw G-lh NS-lh ()
    $width(posedge G, 1.0, 0, notifier);

    // mpw G-hl NS-hl ()
    $width(negedge G, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LARSM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:08:25 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LARSM4N(D, RB, SB, G, Q, QB);
  input D, RB, SB, G;
  output Q, QB;
  reg notifier;

    inv_clr0 SMC_I0(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ));

  `ifdef functional // functional //
    ldlatch_p1 SMC_I2(.q(SMC_IQ), .d(D), .en(G), .clear(RB), .preset(SB));

  `else // functional //
    ldlatch_p1 SMC_I2(.q(SMC_IQ), .d(D), .en(G), .clear(RB), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I6(shcheckGDhl, RB, SB);

    buf SMC_I7(shcheckGRBhl, SB);

    buf SMC_I8(shcheckGSBhl, RB);

    not SMC_I9(shcheckRBSBlh, G);


  specify


    // arc D --> Q
    (D => Q) = (1.0, 1.0);

    // arc D --> QB
    (D => QB) = (1.0, 1.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (1.0, 1.0);

    // arc G --> QB
    (posedge G => ( QB +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl G-hl (RB&SB)
    $setup(negedge D &&& (shcheckGDhl === 1'b1),
        negedge G &&& (shcheckGDhl === 1'b1), 1.0, notifier);

    // setup D-lh G-hl (RB&SB)
    $setup(posedge D &&& (shcheckGDhl === 1'b1),
        negedge G &&& (shcheckGDhl === 1'b1), 1.0, notifier);

    // setup SB-lh RB-lh (!G)
    $setup(posedge SB &&& (shcheckRBSBlh === 1'b1),
        posedge RB &&& (shcheckRBSBlh === 1'b1), 1.0, notifier);

    // hold D-hl G-hl (RB&SB)
    $hold(negedge G &&& (shcheckGDhl === 1'b1),
        negedge D &&& (shcheckGDhl === 1'b1), 1.0, notifier);

    // hold D-lh G-hl (RB&SB)
    $hold(negedge G &&& (shcheckGDhl === 1'b1),
        posedge D &&& (shcheckGDhl === 1'b1), 1.0, notifier);

    // hold SB-lh RB-lh (!G)
    $hold(posedge RB &&& (shcheckRBSBlh === 1'b1),
        posedge SB &&& (shcheckRBSBlh === 1'b1), 1.0, notifier);

    // recovery SB-lh G-hl (RB)
    $recovery(posedge SB &&& (shcheckGSBhl === 1'b1),
        negedge G &&& (shcheckGSBhl === 1'b1), 1.0, notifier);

    // recovery RB-lh G-hl (SB)
    $recovery(posedge RB &&& (shcheckGRBhl === 1'b1),
        negedge G &&& (shcheckGRBhl === 1'b1), 1.0, notifier);

    // removal SB-lh G-hl (RB)
    $hold(negedge G &&& (shcheckGSBhl === 1'b1),
        posedge SB &&& (shcheckGSBhl === 1'b1), 1.0, notifier);

    // removal RB-lh G-hl (SB)
    $hold(negedge G &&& (shcheckGRBhl === 1'b1),
        posedge RB &&& (shcheckGRBhl === 1'b1), 1.0, notifier);

    // mpw G-lh NS-lh ()
    $width(posedge G, 1.0, 0, notifier);

    // mpw G-hl NS-hl ()
    $width(negedge G, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LARSM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:08:25 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LDFQM0N(D, CK, Q);
  input D, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh ()
    $setup(negedge D, posedge CK, 1.0, notifier);

    // setup D-lh CK-lh ()
    $setup(posedge D, posedge CK, 1.0, notifier);

    // hold D-hl CK-lh ()
    $hold(posedge CK, negedge D, 1.0, notifier);

    // hold D-lh CK-lh ()
    $hold(posedge CK, posedge D, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LDFQM0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:08:25 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LDFQM1N(D, CK, Q);
  input D, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh ()
    $setup(negedge D, posedge CK, 1.0, notifier);

    // setup D-lh CK-lh ()
    $setup(posedge D, posedge CK, 1.0, notifier);

    // hold D-hl CK-lh ()
    $hold(posedge CK, negedge D, 1.0, notifier);

    // hold D-lh CK-lh ()
    $hold(posedge CK, posedge D, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LDFQM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:09:09 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LDFQM2N(D, CK, Q);
  input D, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh ()
    $setup(negedge D, posedge CK, 1.0, notifier);

    // setup D-lh CK-lh ()
    $setup(posedge D, posedge CK, 1.0, notifier);

    // hold D-hl CK-lh ()
    $hold(posedge CK, negedge D, 1.0, notifier);

    // hold D-lh CK-lh ()
    $hold(posedge CK, posedge D, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LDFQM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:14:05 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LDFQM4N(D, CK, Q);
  input D, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh ()
    $setup(negedge D, posedge CK, 1.0, notifier);

    // setup D-lh CK-lh ()
    $setup(posedge D, posedge CK, 1.0, notifier);

    // hold D-hl CK-lh ()
    $hold(posedge CK, negedge D, 1.0, notifier);

    // hold D-lh CK-lh ()
    $hold(posedge CK, posedge D, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LDFQM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:14:37 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LDFQRM0N(D, RB, CK, Q);
  input D, RB, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckCKDlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (RB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (RB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 1.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LDFQRM0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:15:39 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LDFQRM1N(D, RB, CK, Q);
  input D, RB, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckCKDlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (RB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (RB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 1.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LDFQRM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:11:02 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LDFQRM2N(D, RB, CK, Q);
  input D, RB, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckCKDlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (RB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (RB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 1.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LDFQRM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:09:20 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LDFQRM4N(D, RB, CK, Q);
  input D, RB, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckCKDlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (RB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (RB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 1.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LDFQRM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:14:10 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LDFQRSM0N(D, RB, SB, CK, Q);
  input D, RB, SB, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //
    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(SB));

  `else // functional //
    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I3(shcheckCKDlh, RB, SB);

    buf SMC_I4(shcheckCKRBlh, SB);

    buf SMC_I5(shcheckCKSBlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);



    // setup SB-lh RB-lh ()
    $setup(posedge SB, posedge RB, 1.0, notifier);

    // setup D-lh CK-lh (RB&SB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (RB&SB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SB-lh RB-lh ()
    $hold(posedge RB, posedge SB, 1.0, notifier);

    // hold D-lh CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh (RB)
    $recovery(posedge SB &&& (shcheckCKSBlh === 1'b1),
        posedge CK &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh (SB)
    $recovery(posedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // removal SB-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSBlh === 1'b1),
        posedge SB &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // removal RB-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        posedge RB &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LDFQRSM0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:13:05 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LDFQRSM1N(D, RB, SB, CK, Q);
  input D, RB, SB, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //
    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(SB));

  `else // functional //
    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I3(shcheckCKDlh, RB, SB);

    buf SMC_I4(shcheckCKRBlh, SB);

    buf SMC_I5(shcheckCKSBlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);



    // setup SB-lh RB-lh ()
    $setup(posedge SB, posedge RB, 1.0, notifier);

    // setup D-lh CK-lh (RB&SB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (RB&SB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SB-lh RB-lh ()
    $hold(posedge RB, posedge SB, 1.0, notifier);

    // hold D-lh CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh (RB)
    $recovery(posedge SB &&& (shcheckCKSBlh === 1'b1),
        posedge CK &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh (SB)
    $recovery(posedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // removal SB-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSBlh === 1'b1),
        posedge SB &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // removal RB-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        posedge RB &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LDFQRSM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:14:28 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LDFQRSM2N(D, RB, SB, CK, Q);
  input D, RB, SB, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //
    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(SB));

  `else // functional //
    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I3(shcheckCKDlh, RB, SB);

    buf SMC_I4(shcheckCKRBlh, SB);

    buf SMC_I5(shcheckCKSBlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);



    // setup SB-lh RB-lh ()
    $setup(posedge SB, posedge RB, 1.0, notifier);

    // setup D-lh CK-lh (RB&SB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (RB&SB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SB-lh RB-lh ()
    $hold(posedge RB, posedge SB, 1.0, notifier);

    // hold D-lh CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh (RB)
    $recovery(posedge SB &&& (shcheckCKSBlh === 1'b1),
        posedge CK &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh (SB)
    $recovery(posedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // removal SB-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSBlh === 1'b1),
        posedge SB &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // removal RB-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        posedge RB &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LDFQRSM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:15:32 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LDFQRSM4N(D, RB, SB, CK, Q);
  input D, RB, SB, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //
    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(SB));

  `else // functional //
    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I3(shcheckCKDlh, RB, SB);

    buf SMC_I4(shcheckCKRBlh, SB);

    buf SMC_I5(shcheckCKSBlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);



    // setup SB-lh RB-lh ()
    $setup(posedge SB, posedge RB, 1.0, notifier);

    // setup D-lh CK-lh (RB&SB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (RB&SB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SB-lh RB-lh ()
    $hold(posedge RB, posedge SB, 1.0, notifier);

    // hold D-lh CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh (RB)
    $recovery(posedge SB &&& (shcheckCKSBlh === 1'b1),
        posedge CK &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh (SB)
    $recovery(posedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // removal SB-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSBlh === 1'b1),
        posedge SB &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // removal RB-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        posedge RB &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LDFQRSM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:08:39 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LDFQSM0N(D, SB, CK, Q);
  input D, SB, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //
    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(SB));

  `else // functional //
    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckCKDlh, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (SB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (SB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 1.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LDFQSM0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:13:45 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LDFQSM1N(D, SB, CK, Q);
  input D, SB, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //
    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(SB));

  `else // functional //
    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckCKDlh, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (SB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (SB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 1.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LDFQSM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:08:39 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LDFQSM2N(D, SB, CK, Q);
  input D, SB, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //
    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(SB));

  `else // functional //
    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckCKDlh, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (SB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (SB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 1.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LDFQSM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:13:18 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LDFQSM4N(D, SB, CK, Q);
  input D, SB, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //
    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(SB));

  `else // functional //
    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckCKDlh, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (SB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (SB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 1.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LDFQSM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:11:39 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LSDFQM0N(D, SD, SE, CK, Q);
  input D, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(shcheckCKDlh, SE);

    buf SMC_I5(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LSDFQM0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:15:46 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LSDFQM1N(D, SD, SE, CK, Q);
  input D, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(shcheckCKDlh, SE);

    buf SMC_I5(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LSDFQM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:08:40 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LSDFQM2N(D, SD, SE, CK, Q);
  input D, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(shcheckCKDlh, SE);

    buf SMC_I5(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LSDFQM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:08:41 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LSDFQM4N(D, SD, SE, CK, Q);
  input D, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(shcheckCKDlh, SE);

    buf SMC_I5(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LSDFQM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:11:09 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LSDFQRM0N(D, RB, SD, SE, CK, Q);
  input D, RB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKDlh, RB, SE_bar);

    and SMC_I6(shcheckCKSDlh, RB, SE);

    buf SMC_I7(shcheckCKSElh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (RB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (RB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (RB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh (RB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (RB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (RB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 1.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LSDFQRM0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:09:25 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LSDFQRM1N(D, RB, SD, SE, CK, Q);
  input D, RB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKDlh, RB, SE_bar);

    and SMC_I6(shcheckCKSDlh, RB, SE);

    buf SMC_I7(shcheckCKSElh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (RB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (RB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (RB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh (RB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (RB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (RB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 1.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LSDFQRM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:14:14 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LSDFQRM2N(D, RB, SD, SE, CK, Q);
  input D, RB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKDlh, RB, SE_bar);

    and SMC_I6(shcheckCKSDlh, RB, SE);

    buf SMC_I7(shcheckCKSElh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (RB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (RB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (RB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh (RB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (RB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (RB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 1.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LSDFQRM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:11:48 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LSDFQRM4N(D, RB, SD, SE, CK, Q);
  input D, RB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKDlh, RB, SE_bar);

    and SMC_I6(shcheckCKSDlh, RB, SE);

    buf SMC_I7(shcheckCKSElh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (RB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (RB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (RB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh (RB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (RB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (RB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 1.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LSDFQRM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:13:57 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LSDFQRSM0N(D, RB, SB, SD, SE, CK, Q);
  input D, RB, SB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(SB));

  `else // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKDlh, RB, SB, SE_bar);

    buf SMC_I6(shcheckCKRBlh, SB);

    buf SMC_I7(shcheckCKSBlh, RB);

    and SMC_I8(shcheckCKSDlh, RB, SB, SE);

    and SMC_I9(shcheckCKSElh, RB, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (RB&SB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (RB&SB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SB-lh RB-lh ()
    $setup(posedge SB, posedge RB, 1.0, notifier);

    // setup SE-hl CK-lh (RB&SB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (RB&SB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (RB&SB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (RB&SB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB&SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB&SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SB-lh RB-lh ()
    $hold(posedge RB, posedge SB, 1.0, notifier);

    // hold SE-hl CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (RB&SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (RB&SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh (SB)
    $recovery(posedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh (RB)
    $recovery(posedge SB &&& (shcheckCKSBlh === 1'b1),
        posedge CK &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // removal RB-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        posedge RB &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // removal SB-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSBlh === 1'b1),
        posedge SB &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LSDFQRSM0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:14:43 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LSDFQRSM1N(D, RB, SB, SD, SE, CK, Q);
  input D, RB, SB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(SB));

  `else // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKDlh, RB, SB, SE_bar);

    buf SMC_I6(shcheckCKRBlh, SB);

    buf SMC_I7(shcheckCKSBlh, RB);

    and SMC_I8(shcheckCKSDlh, RB, SB, SE);

    and SMC_I9(shcheckCKSElh, RB, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (RB&SB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (RB&SB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SB-lh RB-lh ()
    $setup(posedge SB, posedge RB, 1.0, notifier);

    // setup SE-hl CK-lh (RB&SB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (RB&SB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (RB&SB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (RB&SB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB&SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB&SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SB-lh RB-lh ()
    $hold(posedge RB, posedge SB, 1.0, notifier);

    // hold SE-hl CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (RB&SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (RB&SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh (SB)
    $recovery(posedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh (RB)
    $recovery(posedge SB &&& (shcheckCKSBlh === 1'b1),
        posedge CK &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // removal RB-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        posedge RB &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // removal SB-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSBlh === 1'b1),
        posedge SB &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LSDFQRSM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:13:34 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LSDFQRSM2N(D, RB, SB, SD, SE, CK, Q);
  input D, RB, SB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(SB));

  `else // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKDlh, RB, SB, SE_bar);

    buf SMC_I6(shcheckCKRBlh, SB);

    buf SMC_I7(shcheckCKSBlh, RB);

    and SMC_I8(shcheckCKSDlh, RB, SB, SE);

    and SMC_I9(shcheckCKSElh, RB, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (RB&SB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (RB&SB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SB-lh RB-lh ()
    $setup(posedge SB, posedge RB, 1.0, notifier);

    // setup SE-hl CK-lh (RB&SB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (RB&SB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (RB&SB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (RB&SB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB&SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB&SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SB-lh RB-lh ()
    $hold(posedge RB, posedge SB, 1.0, notifier);

    // hold SE-hl CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (RB&SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (RB&SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh (SB)
    $recovery(posedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh (RB)
    $recovery(posedge SB &&& (shcheckCKSBlh === 1'b1),
        posedge CK &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // removal RB-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        posedge RB &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // removal SB-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSBlh === 1'b1),
        posedge SB &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LSDFQRSM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:15:47 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LSDFQRSM4N(D, RB, SB, SD, SE, CK, Q);
  input D, RB, SB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(SB));

  `else // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKDlh, RB, SB, SE_bar);

    buf SMC_I6(shcheckCKRBlh, SB);

    buf SMC_I7(shcheckCKSBlh, RB);

    and SMC_I8(shcheckCKSDlh, RB, SB, SE);

    and SMC_I9(shcheckCKSElh, RB, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (RB&SB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (RB&SB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SB-lh RB-lh ()
    $setup(posedge SB, posedge RB, 1.0, notifier);

    // setup SE-hl CK-lh (RB&SB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (RB&SB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (RB&SB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (RB&SB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB&SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB&SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SB-lh RB-lh ()
    $hold(posedge RB, posedge SB, 1.0, notifier);

    // hold SE-hl CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (RB&SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (RB&SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh (SB)
    $recovery(posedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh (RB)
    $recovery(posedge SB &&& (shcheckCKSBlh === 1'b1),
        posedge CK &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // removal RB-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        posedge RB &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // removal SB-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSBlh === 1'b1),
        posedge SB &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LSDFQRSM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:09:54 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LSDFQSM0N(D, SB, SD, SE, CK, Q);
  input D, SB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(SB));

  `else // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(SB), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKDlh, SB, SE_bar);

    and SMC_I6(shcheckCKSDlh, SB, SE);

    buf SMC_I7(shcheckCKSElh, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (SB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (SB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (SB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh (SB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (SB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 1.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LSDFQSM0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:14:48 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LSDFQSM1N(D, SB, SD, SE, CK, Q);
  input D, SB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(SB));

  `else // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(SB), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKDlh, SB, SE_bar);

    and SMC_I6(shcheckCKSDlh, SB, SE);

    buf SMC_I7(shcheckCKSElh, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (SB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (SB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (SB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh (SB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (SB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 1.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LSDFQSM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:11:39 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LSDFQSM2N(D, SB, SD, SE, CK, Q);
  input D, SB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(SB));

  `else // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(SB), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKDlh, SB, SE_bar);

    and SMC_I6(shcheckCKSDlh, SB, SE);

    buf SMC_I7(shcheckCKSElh, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (SB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (SB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (SB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh (SB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (SB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 1.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LSDFQSM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:15:25 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LSDFQSM4N(D, SB, SD, SE, CK, Q);
  input D, SB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(SB));

  `else // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(SB), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKDlh, SB, SE_bar);

    and SMC_I6(shcheckCKSDlh, SB, SE);

    buf SMC_I7(shcheckCKSElh, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (SB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (SB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (SB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh (SB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (SB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 1.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LSDFQSM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:12:20 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MUX2M0N(A, B, S, Z);
  input A, B, S;
  output Z;

    not SMC_I0(S_bar, S);
    and SMC_I1(OUT0, A, S_bar);
    and SMC_I2(OUT1, B, S);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        (A => Z) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        (B => Z) = (1.0, 1.0);

    // arc S --> Z
     if ( S===1'b1 )
    ( posedge S => ( Z +: S ) ) = (1.0, 1.0);
     if ( S===1'b0 )
    ( negedge S => ( Z +: S ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // MUX2M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 17:23:42 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MUX2M1N(A, B, S, Z);
  input A, B, S;
  output Z;

    not SMC_I0(S_bar, S);
    and SMC_I1(OUT0, A, S_bar);
    and SMC_I2(OUT1, B, S);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        (A => Z) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        (B => Z) = (1.0, 1.0);

    // arc S --> Z
    if (S===1'b1 && S===1'b1 )
    ( posedge S => ( Z +: S ) ) = (1.0, 1.0);
    if (S===1'b0 && S===1'b0 )
    ( negedge S => ( Z +: S ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // MUX2M1N //
`endcelldefine


/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:14:29 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MUX2M2N(A, B, S, Z);
  input A, B, S;
  output Z;

    not SMC_I0(S_bar, S);
    and SMC_I1(OUT0, A, S_bar);
    and SMC_I2(OUT1, B, S);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        (A => Z) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        (B => Z) = (1.0, 1.0);

    // arc S --> Z
     if ( S===1'b1 )
    ( posedge S => ( Z +: S ) ) = (1.0, 1.0);
     if ( S===1'b0 )
    ( negedge S => ( Z +: S ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // MUX2M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:08:58 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MUX2M3N(A, B, S, Z);
  input A, B, S;
  output Z;

    not SMC_I0(S_bar, S);
    and SMC_I1(OUT0, A, S_bar);
    and SMC_I2(OUT1, B, S);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        (A => Z) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        (B => Z) = (1.0, 1.0);

    // arc S --> Z
     if ( S===1'b1 )
    ( posedge S => ( Z +: S ) ) = (1.0, 1.0);
     if ( S===1'b0 )
    ( negedge S => ( Z +: S ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // MUX2M3N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:08:56 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MUX2M4N(A, B, S, Z);
  input A, B, S;
  output Z;

    not SMC_I0(S_bar, S);
    and SMC_I1(OUT0, A, S_bar);
    and SMC_I2(OUT1, B, S);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        (A => Z) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        (B => Z) = (1.0, 1.0);

    // arc S --> Z
     if ( S===1'b1 )
    ( posedge S => ( Z +: S ) ) = (1.0, 1.0);
     if ( S===1'b0 )
    ( negedge S => ( Z +: S ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // MUX2M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:08:58 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MUX2M6N(A, B, S, Z);
  input A, B, S;
  output Z;

    not SMC_I0(S_bar, S);
    and SMC_I1(OUT0, A, S_bar);
    and SMC_I2(OUT1, B, S);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        (A => Z) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        (B => Z) = (1.0, 1.0);

    // arc S --> Z
     if ( S===1'b1 )
    ( posedge S => ( Z +: S ) ) = (1.0, 1.0);
     if ( S===1'b0 )
    ( negedge S => ( Z +: S ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // MUX2M6N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:09:25 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MUX2M8N(A, B, S, Z);
  input A, B, S;
  output Z;

    not SMC_I0(S_bar, S);
    and SMC_I1(OUT0, A, S_bar);
    and SMC_I2(OUT1, B, S);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        (A => Z) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        (B => Z) = (1.0, 1.0);

    // arc S --> Z
     if ( S===1'b1 )
    ( posedge S => ( Z +: S ) ) = (1.0, 1.0);
     if ( S===1'b0 )
    ( negedge S => ( Z +: S ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // MUX2M8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:09:43 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module MUX3M0N ( Z, A, B, C, S0, S1 );
   input A, B, C, S0, S1;
   output Z;
      MUX3M0N_UDP5(Z, A, B, C, S0, S1);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        (A => Z) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        (B => Z) = (1.0, 1.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && S0===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && S0===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && S0===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && S0===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && S0===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && S0===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && S0===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && S0===1'b1) 
        (C => Z) = (1.0, 1.0);
    ifnone
        (C => Z) = (1.0, 1.0);


    // arc S0 --> Z
    if (A===1'b0 && B===1'b1 && C===1'b0 && S1===1'b0)
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && S1===1'b0)
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && S1===1'b0)
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && S1===1'b0)
        (S0 => Z) = (1.0, 1.0);
    ifnone
        (posedge S0 => ( Z +: S0 ) ) = (1.0, 1.0);
        (negedge S0 => ( Z +: S0 ) ) = (1.0, 1.0);


    // arc S1 --> Z
    if (A===1'b0 && B===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    ifnone
        ( posedge S1 => ( Z +: S1 ) ) = (1.0, 1.0);
        ( negedge S1 => ( Z +: S1 ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // MUX3M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:14:07 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module MUX3M1N ( Z, A, B, C, S0, S1 );
   input A, B, C, S0, S1;
   output Z;
      MUX3M0N_UDP5(Z, A, B, C, S0, S1);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        (A => Z) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        (B => Z) = (1.0, 1.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && S0===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && S0===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && S0===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && S0===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && S0===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && S0===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && S0===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && S0===1'b1) 
        (C => Z) = (1.0, 1.0);
    ifnone
        (C => Z) = (1.0, 1.0);

    // arc S0 --> Z
    if (A===1'b0 && B===1'b1 && C===1'b0 && S1===1'b0)
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && S1===1'b0)
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && S1===1'b0)
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && S1===1'b0)
        (S0 => Z) = (1.0, 1.0);
    ifnone
        (posedge S0 => ( Z +: S0 ) ) = (1.0, 1.0);
        (negedge S0 => ( Z +: S0 ) ) = (1.0, 1.0);

    // arc S1 --> Z
    if (A===1'b0 && B===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    ifnone
        ( posedge S1 => ( Z +: S1 ) ) = (1.0, 1.0);
        ( negedge S1 => ( Z +: S1 ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // MUX3M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:17:38 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module MUX3M2N ( Z, A, B, C, S0, S1 );
   input A, B, C, S0, S1;
   output Z;
      MUX3M0N_UDP5(Z, A, B, C, S0, S1);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        (A => Z) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        (B => Z) = (1.0, 1.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && S0===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && S0===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && S0===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && S0===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && S0===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && S0===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && S0===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && S0===1'b1) 
        (C => Z) = (1.0, 1.0);
    ifnone
        (C => Z) = (1.0, 1.0);


    // arc S0 --> Z
    if (A===1'b0 && B===1'b1 && C===1'b0 && S1===1'b0)
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && S1===1'b0)
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && S1===1'b0)
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && S1===1'b0)
        (S0 => Z) = (1.0, 1.0);
    ifnone
        (posedge S0 => ( Z +: S0 ) ) = (1.0, 1.0);
        (negedge S0 => ( Z +: S0 ) ) = (1.0, 1.0);

    // arc S1 --> Z
    if (A===1'b0 && B===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    ifnone
        ( posedge S1 => ( Z +: S1 ) ) = (1.0, 1.0);
        ( negedge S1 => ( Z +: S1 ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // MUX3M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:13:20 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module MUX3M4N ( Z, A, B, C, S0, S1 );
   input A, B, C, S0, S1;
   output Z;
      MUX3M0N_UDP5(Z, A, B, C, S0, S1);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        (A => Z) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        (B => Z) = (1.0, 1.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && S0===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && S0===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && S0===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && S0===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && S0===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && S0===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && S0===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && S0===1'b1) 
        (C => Z) = (1.0, 1.0);
    ifnone
        (C => Z) = (1.0, 1.0);

    // arc S0 --> Z
    if (A===1'b0 && B===1'b1 && C===1'b0 && S1===1'b0)
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && S1===1'b0)
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && S1===1'b0)
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && S1===1'b0)
        (S0 => Z) = (1.0, 1.0);
    ifnone
        (posedge S0 => ( Z +: S0 ) ) = (1.0, 1.0);
        (negedge S0 => ( Z +: S0 ) ) = (1.0, 1.0);


    // arc S1 --> Z
    if (A===1'b0 && B===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    ifnone
        ( posedge S1 => ( Z +: S1 ) ) = (1.0, 1.0);
        ( negedge S1 => ( Z +: S1 ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // MUX3M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:11:55 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module MUX4M0N ( Z, A, B, C, D, S0, S1 );
   input A, B, C, D, S0, S1;
   output Z;
      MUX4M0N_UDP6(Z, A, B, C, D, S0, S1);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0 && D===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b0 && C===1'b0 && D===1'b1) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1 && D===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1 && D===1'b1) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0 && D===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0 && D===1'b1) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1 && D===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1 && D===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        (A => Z) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0 && D===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b0 && C===1'b0 && D===1'b1) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1 && D===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1 && D===1'b1) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0 && D===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0 && D===1'b1) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1 && D===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1 && D===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        (B => Z) = (1.0, 1.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && D===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && D===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && D===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && D===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && D===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && D===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && D===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && D===1'b1) 
        (C => Z) = (1.0, 1.0);
    ifnone
        (C => Z) = (1.0, 1.0);

    // arc D --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b1) 
        (D => Z) = (1.0, 1.0);
    ifnone
        (D => Z) = (1.0, 1.0);

    // arc S0 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    ifnone
        ( posedge S0 => ( Z +: S0 ) ) = (1.0, 1.0);
        ( negedge S0 => ( Z +: S0 ) ) = (1.0, 1.0);

    // arc S1 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    ifnone
        ( posedge S1 => ( Z +: S1 ) ) = (1.0, 1.0);
        ( negedge S1 => ( Z +: S1 ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // MUX4M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:14:48 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module MUX4M1N ( Z, A, B, C, D, S0, S1 );
   input A, B, C, D, S0, S1;
   output Z;
      MUX4M0N_UDP6(Z, A, B, C, D, S0, S1);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0 && D===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b0 && C===1'b0 && D===1'b1) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1 && D===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1 && D===1'b1) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0 && D===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0 && D===1'b1) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1 && D===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1 && D===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        (A => Z) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0 && D===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b0 && C===1'b0 && D===1'b1) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1 && D===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1 && D===1'b1) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0 && D===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0 && D===1'b1) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1 && D===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1 && D===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        (B => Z) = (1.0, 1.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && D===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && D===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && D===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && D===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && D===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && D===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && D===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && D===1'b1) 
        (C => Z) = (1.0, 1.0);
    ifnone
        (C => Z) = (1.0, 1.0);

    // arc D --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b1) 
        (D => Z) = (1.0, 1.0);
    ifnone
        (D => Z) = (1.0, 1.0);

    // arc S0 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    ifnone
        ( posedge S0 => ( Z +: S0 ) ) = (1.0, 1.0);
        ( negedge S0 => ( Z +: S0 ) ) = (1.0, 1.0);

    // arc S1 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    ifnone
        ( posedge S1 => ( Z +: S1 ) ) = (1.0, 1.0);
        ( negedge S1 => ( Z +: S1 ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // MUX4M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:11:20 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module MUX4M2N ( Z, A, B, C, D, S0, S1 );
   input A, B, C, D, S0, S1;
   output Z;
      MUX4M0N_UDP6(Z, A, B, C, D, S0, S1);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0 && D===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b0 && C===1'b0 && D===1'b1) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1 && D===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1 && D===1'b1) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0 && D===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0 && D===1'b1) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1 && D===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1 && D===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        (A => Z) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0 && D===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b0 && C===1'b0 && D===1'b1) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1 && D===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1 && D===1'b1) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0 && D===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0 && D===1'b1) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1 && D===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1 && D===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        (B => Z) = (1.0, 1.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && D===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && D===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && D===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && D===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && D===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && D===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && D===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && D===1'b1) 
        (C => Z) = (1.0, 1.0);
    ifnone
        (C => Z) = (1.0, 1.0);

    // arc D --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b1) 
        (D => Z) = (1.0, 1.0);
    ifnone
        (D => Z) = (1.0, 1.0);

    // arc S0 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    ifnone
        ( posedge S0 => ( Z +: S0 ) ) = (1.0, 1.0);
        ( negedge S0 => ( Z +: S0 ) ) = (1.0, 1.0);

    // arc S1 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    ifnone
        ( posedge S1 => ( Z +: S1 ) ) = (1.0, 1.0);
        ( negedge S1 => ( Z +: S1 ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // MUX4M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:16:18 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module MUX4M4N ( Z, A, B, C, D, S0, S1 );
   input A, B, C, D, S0, S1;
   output Z;
      MUX4M0N_UDP6(Z, A, B, C, D, S0, S1);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0 && D===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b0 && C===1'b0 && D===1'b1) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1 && D===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1 && D===1'b1) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0 && D===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0 && D===1'b1) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1 && D===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1 && D===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        (A => Z) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0 && D===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b0 && C===1'b0 && D===1'b1) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1 && D===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1 && D===1'b1) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0 && D===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0 && D===1'b1) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1 && D===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1 && D===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        (B => Z) = (1.0, 1.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && D===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && D===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && D===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && D===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && D===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && D===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && D===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && D===1'b1) 
        (C => Z) = (1.0, 1.0);
    ifnone
        (C => Z) = (1.0, 1.0);

    // arc D --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b1) 
        (D => Z) = (1.0, 1.0);
    ifnone
        (D => Z) = (1.0, 1.0);

    // arc S0 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    ifnone
        ( posedge S0 => ( Z +: S0 ) ) = (1.0, 1.0);
        ( negedge S0 => ( Z +: S0 ) ) = (1.0, 1.0);

    // arc S1 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    ifnone
        ( posedge S1 => ( Z +: S1 ) ) = (1.0, 1.0);
        ( negedge S1 => ( Z +: S1 ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // MUX4M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:16:35 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MXB2DM0N(A, B, S, Z);
  input A, B, S;
  output Z;

    not SMC_I0(A_bar, A);
    not SMC_I1(S_bar, S);
    and SMC_I2(OUT0, A_bar, S_bar);
    not SMC_I3(B_bar, B);
    and SMC_I4(OUT1, B_bar, S);
    or SMC_I5(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        (A => Z) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        (B => Z) = (1.0, 1.0);

    // arc S --> Z
     if ( S===1'b1 )
    ( posedge S => ( Z +: S ) ) = (1.0, 1.0);
     if ( S===1'b0 )
    ( negedge S => ( Z +: S ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // MXB2DM0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:13:39 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MXB2DM1N(A, B, S, Z);
  input A, B, S;
  output Z;

    not SMC_I0(A_bar, A);
    not SMC_I1(S_bar, S);
    and SMC_I2(OUT0, A_bar, S_bar);
    not SMC_I3(B_bar, B);
    and SMC_I4(OUT1, B_bar, S);
    or SMC_I5(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        (A => Z) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        (B => Z) = (1.0, 1.0);

    // arc S --> Z
     if ( S===1'b1 )
    ( posedge S => ( Z +: S ) ) = (1.0, 1.0);
     if ( S===1'b0 )
    ( negedge S => ( Z +: S ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // MXB2DM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:18:32 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MXB2DM2N(A, B, S, Z);
  input A, B, S;
  output Z;

    not SMC_I0(A_bar, A);
    not SMC_I1(S_bar, S);
    and SMC_I2(OUT0, A_bar, S_bar);
    not SMC_I3(B_bar, B);
    and SMC_I4(OUT1, B_bar, S);
    or SMC_I5(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        (A => Z) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        (B => Z) = (1.0, 1.0);

    // arc S --> Z
     if ( S===1'b1 )
    ( posedge S => ( Z +: S ) ) = (1.0, 1.0);
     if ( S===1'b0 )
    ( negedge S => ( Z +: S ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // MXB2DM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:11:34 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MXB2DM4N(A, B, S, Z);
  input A, B, S;
  output Z;

    not SMC_I0(A_bar, A);
    not SMC_I1(S_bar, S);
    and SMC_I2(OUT0, A_bar, S_bar);
    not SMC_I3(B_bar, B);
    and SMC_I4(OUT1, B_bar, S);
    or SMC_I5(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        (A => Z) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        (B => Z) = (1.0, 1.0);

    // arc S --> Z
     if ( S===1'b1 )
    ( posedge S => ( Z +: S ) ) = (1.0, 1.0);
     if ( S===1'b0 )
    ( negedge S => ( Z +: S ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // MXB2DM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:11:28 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MXB2M0N(A, B, S, Z);
  input A, B, S;
  output Z;

    not SMC_I0(A_bar, A);
    not SMC_I1(S_bar, S);
    and SMC_I2(OUT0, A_bar, S_bar);
    not SMC_I3(B_bar, B);
    and SMC_I4(OUT1, B_bar, S);
    or SMC_I5(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        (A => Z) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        (B => Z) = (1.0, 1.0);

    // arc S --> Z
     if ( S===1'b1 )
    ( posedge S => ( Z +: S ) ) = (1.0, 1.0);
     if ( S===1'b0 )
    ( negedge S => ( Z +: S ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // MXB2M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:11:37 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MXB2M1N(A, B, S, Z);
  input A, B, S;
  output Z;

    not SMC_I0(A_bar, A);
    not SMC_I1(S_bar, S);
    and SMC_I2(OUT0, A_bar, S_bar);
    not SMC_I3(B_bar, B);
    and SMC_I4(OUT1, B_bar, S);
    or SMC_I5(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        (A => Z) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        (B => Z) = (1.0, 1.0);

    // arc S --> Z
     if ( S===1'b1 )
    ( posedge S => ( Z +: S ) ) = (1.0, 1.0);
     if ( S===1'b0 )
    ( negedge S => ( Z +: S ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // MXB2M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:11:35 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MXB2M2N(A, B, S, Z);
  input A, B, S;
  output Z;

    not SMC_I0(A_bar, A);
    not SMC_I1(S_bar, S);
    and SMC_I2(OUT0, A_bar, S_bar);
    not SMC_I3(B_bar, B);
    and SMC_I4(OUT1, B_bar, S);
    or SMC_I5(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        (A => Z) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        (B => Z) = (1.0, 1.0);

    // arc S --> Z
     if ( S===1'b1 )
    ( posedge S => ( Z +: S ) ) = (1.0, 1.0);
     if ( S===1'b0 )
    ( negedge S => ( Z +: S ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // MXB2M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:14:29 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MXB2M3N(A, B, S, Z);
  input A, B, S;
  output Z;

    not SMC_I0(A_bar, A);
    not SMC_I1(S_bar, S);
    and SMC_I2(OUT0, A_bar, S_bar);
    not SMC_I3(B_bar, B);
    and SMC_I4(OUT1, B_bar, S);
    or SMC_I5(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        (A => Z) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        (B => Z) = (1.0, 1.0);

    // arc S --> Z
     if ( S===1'b1 )
    ( posedge S => ( Z +: S ) ) = (1.0, 1.0);
     if ( S===1'b0 )
    ( negedge S => ( Z +: S ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // MXB2M3N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:11:35 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MXB2M4N(A, B, S, Z);
  input A, B, S;
  output Z;

    not SMC_I0(A_bar, A);
    not SMC_I1(S_bar, S);
    and SMC_I2(OUT0, A_bar, S_bar);
    not SMC_I3(B_bar, B);
    and SMC_I4(OUT1, B_bar, S);
    or SMC_I5(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        (A => Z) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        (B => Z) = (1.0, 1.0);

    // arc S --> Z
     if ( S===1'b1 )
    ( posedge S => ( Z +: S ) ) = (1.0, 1.0);
     if ( S===1'b0 )
    ( negedge S => ( Z +: S ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // MXB2M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:14:42 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MXB2M6N(A, B, S, Z);
  input A, B, S;
  output Z;

    not SMC_I0(A_bar, A);
    not SMC_I1(S_bar, S);
    and SMC_I2(OUT0, A_bar, S_bar);
    not SMC_I3(B_bar, B);
    and SMC_I4(OUT1, B_bar, S);
    or SMC_I5(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        (A => Z) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        (B => Z) = (1.0, 1.0);

    // arc S --> Z
     if ( S===1'b1 )
    ( posedge S => ( Z +: S ) ) = (1.0, 1.0);
     if ( S===1'b0 )
    ( negedge S => ( Z +: S ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // MXB2M6N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:15:12 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MXB2M8N(A, B, S, Z);
  input A, B, S;
  output Z;

    not SMC_I0(A_bar, A);
    not SMC_I1(S_bar, S);
    and SMC_I2(OUT0, A_bar, S_bar);
    not SMC_I3(B_bar, B);
    and SMC_I4(OUT1, B_bar, S);
    or SMC_I5(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        (A => Z) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        (B => Z) = (1.0, 1.0);

    // arc S --> Z
     if ( S===1'b1 )
    ( posedge S => ( Z +: S ) ) = (1.0, 1.0);
     if ( S===1'b0 )
    ( negedge S => ( Z +: S ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // MXB2M8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:13:50 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module MXB3M0N ( Z, A, B, C, S0, S1 );
   input A, B, C, S0, S1;
   output Z;
      MXB3M0N_UDP5(Z, A, B, C, S0, S1);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        (A => Z) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        (B => Z) = (1.0, 1.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && S0===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && S0===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && S0===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && S0===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && S0===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && S0===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && S0===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && S0===1'b1) 
        (C => Z) = (1.0, 1.0);
    ifnone
        (C => Z) = (1.0, 1.0);

    // arc S0 --> Z
    if (A===1'b0 && B===1'b1 && C===1'b0 && S1===1'b0)
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && S1===1'b0)
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && S1===1'b0)
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && S1===1'b0)
        (S0 => Z) = (1.0, 1.0);
    ifnone
        (posedge S0 => ( Z +: S0 ) ) = (1.0, 1.0);
        (negedge S0 => ( Z +: S0 ) ) = (1.0, 1.0);


    // arc S1 --> Z
    if (A===1'b0 && B===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    ifnone
        ( posedge S1 => ( Z +: S1 ) ) = (1.0, 1.0);
        ( negedge S1 => ( Z +: S1 ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // MXB3M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:11:38 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module MXB3M1N ( Z, A, B, C, S0, S1 );
   input A, B, C, S0, S1;
   output Z;
      MXB3M0N_UDP5(Z, A, B, C, S0, S1);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        (A => Z) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        (B => Z) = (1.0, 1.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && S0===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && S0===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && S0===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && S0===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && S0===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && S0===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && S0===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && S0===1'b1) 
        (C => Z) = (1.0, 1.0);
    ifnone
        (C => Z) = (1.0, 1.0);


    // arc S0 --> Z
    if (A===1'b0 && B===1'b1 && C===1'b0 && S1===1'b0)
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && S1===1'b0)
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && S1===1'b0)
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && S1===1'b0)
        (S0 => Z) = (1.0, 1.0);
    ifnone
        (posedge S0 => ( Z +: S0 ) ) = (1.0, 1.0);
        (negedge S0 => ( Z +: S0 ) ) = (1.0, 1.0);

    // arc S1 --> Z
    if (A===1'b0 && B===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    ifnone
        ( posedge S1 => ( Z +: S1 ) ) = (1.0, 1.0);
        ( negedge S1 => ( Z +: S1 ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // MXB3M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:16:16 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module MXB3M2N ( Z, A, B, C, S0, S1 );
   input A, B, C, S0, S1;
   output Z;
      MXB3M0N_UDP5(Z, A, B, C, S0, S1);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        (A => Z) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        (B => Z) = (1.0, 1.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && S0===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && S0===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && S0===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && S0===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && S0===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && S0===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && S0===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && S0===1'b1) 
        (C => Z) = (1.0, 1.0);
    ifnone
        (C => Z) = (1.0, 1.0);

    // arc S0 --> Z
    if (A===1'b0 && B===1'b1 && C===1'b0 && S1===1'b0)
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && S1===1'b0)
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && S1===1'b0)
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && S1===1'b0)
        (S0 => Z) = (1.0, 1.0);
    ifnone
        (posedge S0 => ( Z +: S0 ) ) = (1.0, 1.0);
        (negedge S0 => ( Z +: S0 ) ) = (1.0, 1.0);

    // arc S1 --> Z
    if (A===1'b0 && B===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    ifnone
        ( posedge S1 => ( Z +: S1 ) ) = (1.0, 1.0);
        ( negedge S1 => ( Z +: S1 ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // MXB3M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:12:29 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module MXB3M4N ( Z, A, B, C, S0, S1 );
   input A, B, C, S0, S1;
   output Z;
      MXB3M0N_UDP5(Z, A, B, C, S0, S1);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        (A => Z) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        (B => Z) = (1.0, 1.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && S0===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && S0===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && S0===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && S0===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && S0===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && S0===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && S0===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && S0===1'b1) 
        (C => Z) = (1.0, 1.0);
    ifnone
        (C => Z) = (1.0, 1.0);

    // arc S0 --> Z
    if (A===1'b0 && B===1'b1 && C===1'b0 && S1===1'b0)
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && S1===1'b0)
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && S1===1'b0)
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && S1===1'b0)
        (S0 => Z) = (1.0, 1.0);
    ifnone
        (posedge S0 => ( Z +: S0 ) ) = (1.0, 1.0);
        (negedge S0 => ( Z +: S0 ) ) = (1.0, 1.0);

    // arc S1 --> Z
    if (A===1'b0 && B===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    ifnone
        ( posedge S1 => ( Z +: S1 ) ) = (1.0, 1.0);
        ( negedge S1 => ( Z +: S1 ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // MXB3M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:12:49 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module MXB4M0N ( Z, A, B, C, D, S0, S1 );
   input A, B, C, D, S0, S1;
   output Z;
      MXB4M0N_UDP6(Z, A, B, C, D, S0, S1);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0 && D===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b0 && C===1'b0 && D===1'b1) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1 && D===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1 && D===1'b1) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0 && D===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0 && D===1'b1) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1 && D===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1 && D===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        (A => Z) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0 && D===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b0 && C===1'b0 && D===1'b1) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1 && D===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1 && D===1'b1) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0 && D===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0 && D===1'b1) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1 && D===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1 && D===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        (B => Z) = (1.0, 1.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && D===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && D===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && D===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && D===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && D===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && D===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && D===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && D===1'b1) 
        (C => Z) = (1.0, 1.0);
    ifnone
        (C => Z) = (1.0, 1.0);

    // arc D --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b1) 
        (D => Z) = (1.0, 1.0);
    ifnone
        (D => Z) = (1.0, 1.0);

    // arc S0 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    ifnone
        ( posedge S0 => ( Z +: S0 ) ) = (1.0, 1.0);
        ( negedge S0 => ( Z +: S0 ) ) = (1.0, 1.0);

    // arc S1 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    ifnone
        ( posedge S1 => ( Z +: S1 ) ) = (1.0, 1.0);
        ( negedge S1 => ( Z +: S1 ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // MXB4M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:16:46 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module MXB4M1N ( Z, A, B, C, D, S0, S1 );
   input A, B, C, D, S0, S1;
   output Z;
      MXB4M0N_UDP6(Z, A, B, C, D, S0, S1);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0 && D===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b0 && C===1'b0 && D===1'b1) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1 && D===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1 && D===1'b1) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0 && D===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0 && D===1'b1) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1 && D===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1 && D===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        (A => Z) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0 && D===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b0 && C===1'b0 && D===1'b1) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1 && D===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1 && D===1'b1) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0 && D===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0 && D===1'b1) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1 && D===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1 && D===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        (B => Z) = (1.0, 1.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && D===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && D===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && D===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && D===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && D===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && D===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && D===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && D===1'b1) 
        (C => Z) = (1.0, 1.0);
    ifnone
        (C => Z) = (1.0, 1.0);

    // arc D --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b1) 
        (D => Z) = (1.0, 1.0);
    ifnone
        (D => Z) = (1.0, 1.0);

    // arc S0 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    ifnone
        ( posedge S0 => ( Z +: S0 ) ) = (1.0, 1.0);
        ( negedge S0 => ( Z +: S0 ) ) = (1.0, 1.0);

    // arc S1 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    ifnone
        ( posedge S1 => ( Z +: S1 ) ) = (1.0, 1.0);
        ( negedge S1 => ( Z +: S1 ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // MXB4M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:12:43 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module MXB4M2N ( Z, A, B, C, D, S0, S1 );
   input A, B, C, D, S0, S1;
   output Z;
      MXB4M0N_UDP6(Z, A, B, C, D, S0, S1);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0 && D===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b0 && C===1'b0 && D===1'b1) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1 && D===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1 && D===1'b1) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0 && D===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0 && D===1'b1) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1 && D===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1 && D===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        (A => Z) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0 && D===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b0 && C===1'b0 && D===1'b1) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1 && D===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1 && D===1'b1) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0 && D===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0 && D===1'b1) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1 && D===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1 && D===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        (B => Z) = (1.0, 1.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && D===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && D===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && D===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && D===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && D===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && D===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && D===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && D===1'b1) 
        (C => Z) = (1.0, 1.0);
    ifnone
        (C => Z) = (1.0, 1.0);

    // arc D --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b1) 
        (D => Z) = (1.0, 1.0);
    ifnone
        (D => Z) = (1.0, 1.0);

    // arc S0 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    ifnone
        ( posedge S0 => ( Z +: S0 ) ) = (1.0, 1.0);
        ( negedge S0 => ( Z +: S0 ) ) = (1.0, 1.0);

    // arc S1 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    ifnone
        ( posedge S1 => ( Z +: S1 ) ) = (1.0, 1.0);
        ( negedge S1 => ( Z +: S1 ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // MXB4M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:11:49 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module MXB4M4N ( Z, A, B, C, D, S0, S1 );
   input A, B, C, D, S0, S1;
   output Z;
      MXB4M0N_UDP6(Z, A, B, C, D, S0, S1);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0 && D===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b0 && C===1'b0 && D===1'b1) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1 && D===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1 && D===1'b1) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0 && D===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0 && D===1'b1) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1 && D===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1 && D===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        (A => Z) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0 && D===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b0 && C===1'b0 && D===1'b1) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1 && D===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1 && D===1'b1) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0 && D===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0 && D===1'b1) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1 && D===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1 && D===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        (B => Z) = (1.0, 1.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && D===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && D===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && D===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && D===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && D===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && D===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && D===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && D===1'b1) 
        (C => Z) = (1.0, 1.0);
    ifnone
        (C => Z) = (1.0, 1.0);

    // arc D --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0) 
        (D => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b1) 
        (D => Z) = (1.0, 1.0);
    ifnone
        (D => Z) = (1.0, 1.0);

    // arc S0 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S1===1'b0) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1) 
        (S0 => Z) = (1.0, 1.0);
    ifnone
        ( posedge S0 => ( Z +: S0 ) ) = (1.0, 1.0);
        ( negedge S0 => ( Z +: S0 ) ) = (1.0, 1.0);

    // arc S1 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0) 
        (S1 => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1) 
        (S1 => Z) = (1.0, 1.0);
    ifnone
        ( posedge S1 => ( Z +: S1 ) ) = (1.0, 1.0);
        ( negedge S1 => ( Z +: S1 ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // MXB4M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:12:24 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND2B1M0N(B, NA, Z);
  input B, NA;
  output Z;

    not SMC_I0(NA_bar, NA);
    nand SMC_I1(Z, B, NA_bar);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc NA --> Z
    (NA => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ND2B1M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:14:57 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND2B1M1N(B, NA, Z);
  input B, NA;
  output Z;

    not SMC_I0(NA_bar, NA);
    nand SMC_I1(Z, B, NA_bar);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc NA --> Z
    (NA => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ND2B1M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:10:09 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND2B1M2N(B, NA, Z);
  input B, NA;
  output Z;

    not SMC_I0(NA_bar, NA);
    nand SMC_I1(Z, B, NA_bar);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc NA --> Z
    (NA => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ND2B1M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:11:50 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND2B1M4N(B, NA, Z);
  input B, NA;
  output Z;

    not SMC_I0(NA_bar, NA);
    nand SMC_I1(Z, B, NA_bar);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc NA --> Z
    (NA => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ND2B1M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:15:27 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND2B1M8N(B, NA, Z);
  input B, NA;
  output Z;

    not SMC_I0(NA_bar, NA);
    nand SMC_I1(Z, B, NA_bar);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc NA --> Z
    (NA => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ND2B1M8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:17:30 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND2M0N(A, B, Z);
  input A, B;
  output Z;

    nand SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ND2M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:15:52 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND2M1N(A, B, Z);
  input A, B;
  output Z;

    nand SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ND2M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:18:26 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND2M2N(A, B, Z);
  input A, B;
  output Z;

    nand SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ND2M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:14:32 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND2M3N(A, B, Z);
  input A, B;
  output Z;

    nand SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ND2M3N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:10:11 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND2M4N(A, B, Z);
  input A, B;
  output Z;

    nand SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ND2M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:11:52 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND2M5N(A, B, Z);
  input A, B;
  output Z;

    nand SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ND2M5N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:15:41 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND2M6N(A, B, Z);
  input A, B;
  output Z;

    nand SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ND2M6N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:14:46 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND2M8N(A, B, Z);
  input A, B;
  output Z;

    nand SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ND2M8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:10:24 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module ND3B1M0N ( Z, B, C, NA );
   input B, C, NA;
   output Z;
      ND3B1M0N_UDP3(Z, B, C, NA);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc NA --> Z
    (NA => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ND3B1M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:15:12 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module ND3B1M1N ( Z, B, C, NA );
   input B, C, NA;
   output Z;
      ND3B1M0N_UDP3(Z, B, C, NA);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc NA --> Z
    (NA => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ND3B1M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:12:05 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module ND3B1M2N ( Z, B, C, NA );
   input B, C, NA;
   output Z;
      ND3B1M0N_UDP3(Z, B, C, NA);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc NA --> Z
    (NA => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ND3B1M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:17:36 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module ND3B1M4N ( Z, B, C, NA );
   input B, C, NA;
   output Z;
      ND3B1M0N_UDP3(Z, B, C, NA);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc NA --> Z
    (NA => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ND3B1M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:18:56 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module ND3M0N ( Z, A, B, C );
   input A, B, C;
   output Z;
      ND3M0N_UDP3(Z, A, B, C);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ND3M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:15:27 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module ND3M1N ( Z, A, B, C );
   input A, B, C;
   output Z;
      ND3M0N_UDP3(Z, A, B, C);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ND3M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:15:01 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module ND3M2N ( Z, A, B, C );
   input A, B, C;
   output Z;
      ND3M0N_UDP3(Z, A, B, C);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ND3M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:10:39 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module ND3M3N ( Z, A, B, C );
   input A, B, C;
   output Z;
      ND3M0N_UDP3(Z, A, B, C);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ND3M3N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:12:20 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module ND3M4N ( Z, A, B, C );
   input A, B, C;
   output Z;
      ND3M0N_UDP3(Z, A, B, C);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ND3M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:15:57 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module ND3M6N ( Z, A, B, C );
   input A, B, C;
   output Z;
      ND3M0N_UDP3(Z, A, B, C);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ND3M6N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:20:04 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module ND3M8N ( Z, A, B, C );
   input A, B, C;
   output Z;
      ND3M0N_UDP3(Z, A, B, C);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ND3M8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:13:09 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module ND4B1M0N ( Z, B, C, D, NA );
   input B, C, D, NA;
   output Z;
      ND4B1M0N_UDP4(Z, B, C, D, NA);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc D --> Z
    (D => Z) = (1.0, 1.0);

    // arc NA --> Z
    (NA => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ND4B1M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:17:39 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module ND4B1M1N ( Z, B, C, D, NA );
   input B, C, D, NA;
   output Z;
      ND4B1M0N_UDP4(Z, B, C, D, NA);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc D --> Z
    (D => Z) = (1.0, 1.0);

    // arc NA --> Z
    (NA => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ND4B1M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:16:03 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module ND4B1M2N ( Z, B, C, D, NA );
   input B, C, D, NA;
   output Z;
      ND4B1M0N_UDP4(Z, B, C, D, NA);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc D --> Z
    (D => Z) = (1.0, 1.0);

    // arc NA --> Z
    (NA => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ND4B1M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:18:39 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module ND4B1M4N ( Z, B, C, D, NA );
   input B, C, D, NA;
   output Z;
      ND4B1M0N_UDP4(Z, B, C, D, NA);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc D --> Z
    (D => Z) = (1.0, 1.0);

    // arc NA --> Z
    (NA => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ND4B1M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:13:58 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module ND4B2M0N ( Z, C, D, NA, NB );
   input C, D, NA, NB;
   output Z;
      ND4B2M0N_UDP4(Z, C, D, NA, NB);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc D --> Z
    (D => Z) = (1.0, 1.0);

    // arc NA --> Z
    (NA => Z) = (1.0, 1.0);

    // arc NB --> Z
    (NB => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ND4B2M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:18:23 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module ND4B2M1N ( Z, C, D, NA, NB );
   input C, D, NA, NB;
   output Z;
      ND4B2M0N_UDP4(Z, C, D, NA, NB);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc D --> Z
    (D => Z) = (1.0, 1.0);

    // arc NA --> Z
    (NA => Z) = (1.0, 1.0);

    // arc NB --> Z
    (NB => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ND4B2M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:15:45 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module ND4B2M2N ( Z, C, D, NA, NB );
   input C, D, NA, NB;
   output Z;
      ND4B2M0N_UDP4(Z, C, D, NA, NB);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc D --> Z
    (D => Z) = (1.0, 1.0);

    // arc NA --> Z
    (NA => Z) = (1.0, 1.0);

    // arc NB --> Z
    (NB => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ND4B2M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:19:30 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module ND4B2M4N ( Z, C, D, NA, NB );
   input C, D, NA, NB;
   output Z;
      ND4B2M0N_UDP4(Z, C, D, NA, NB);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc D --> Z
    (D => Z) = (1.0, 1.0);

    // arc NA --> Z
    (NA => Z) = (1.0, 1.0);

    // arc NB --> Z
    (NB => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ND4B2M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:20:28 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module ND4M0N ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;
      ND4M0N_UDP4(Z, A, B, C, D);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc D --> Z
    (D => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ND4M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:18:04 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module ND4M1N ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;
      ND4M0N_UDP4(Z, A, B, C, D);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc D --> Z
    (D => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ND4M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:10:58 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module ND4M2N ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;
      ND4M0N_UDP4(Z, A, B, C, D);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc D --> Z
    (D => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ND4M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:15:45 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module ND4M4N ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;
      ND4M0N_UDP4(Z, A, B, C, D);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc D --> Z
    (D => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ND4M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:15:20 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module ND4M6N ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;
      ND4M0N_UDP4(Z, A, B, C, D);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc D --> Z
    (D => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ND4M6N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:16:16 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module ND4M8N ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;
      ND4M0N_UDP4(Z, A, B, C, D);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc D --> Z
    (D => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ND4M8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:12:39 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR2B1M0N(B, NA, Z);
  input B, NA;
  output Z;

    not SMC_I0(B_bar, B);
    and SMC_I1(Z, B_bar, NA);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc NA --> Z
    (NA => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // NR2B1M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:13:05 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR2B1M1N(B, NA, Z);
  input B, NA;
  output Z;

    not SMC_I0(B_bar, B);
    and SMC_I1(Z, B_bar, NA);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc NA --> Z
    (NA => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // NR2B1M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:16:41 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR2B1M2N(B, NA, Z);
  input B, NA;
  output Z;

    not SMC_I0(B_bar, B);
    and SMC_I1(Z, B_bar, NA);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc NA --> Z
    (NA => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // NR2B1M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:15:46 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR2B1M4N(B, NA, Z);
  input B, NA;
  output Z;

    not SMC_I0(B_bar, B);
    and SMC_I1(Z, B_bar, NA);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc NA --> Z
    (NA => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // NR2B1M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:13:40 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR2B1M8N(B, NA, Z);
  input B, NA;
  output Z;

    not SMC_I0(B_bar, B);
    and SMC_I1(Z, B_bar, NA);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc NA --> Z
    (NA => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // NR2B1M8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:19:04 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR2M0N(A, B, Z);
  input A, B;
  output Z;

    not SMC_I0(A_bar, A);
    not SMC_I1(B_bar, B);
    and SMC_I2(Z, A_bar, B_bar);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // NR2M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:11:24 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR2M1N(A, B, Z);
  input A, B;
  output Z;

    not SMC_I0(A_bar, A);
    not SMC_I1(B_bar, B);
    and SMC_I2(Z, A_bar, B_bar);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // NR2M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:13:05 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR2M2N(A, B, Z);
  input A, B;
  output Z;

    not SMC_I0(A_bar, A);
    not SMC_I1(B_bar, B);
    and SMC_I2(Z, A_bar, B_bar);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // NR2M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:13:20 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR2M3N(A, B, Z);
  input A, B;
  output Z;

    not SMC_I0(A_bar, A);
    not SMC_I1(B_bar, B);
    and SMC_I2(Z, A_bar, B_bar);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // NR2M3N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:16:56 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR2M4N(A, B, Z);
  input A, B;
  output Z;

    not SMC_I0(A_bar, A);
    not SMC_I1(B_bar, B);
    and SMC_I2(Z, A_bar, B_bar);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // NR2M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:16:01 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR2M5N(A, B, Z);
  input A, B;
  output Z;

    not SMC_I0(A_bar, A);
    not SMC_I1(B_bar, B);
    and SMC_I2(Z, A_bar, B_bar);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // NR2M5N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:13:55 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR2M6N(A, B, Z);
  input A, B;
  output Z;

    not SMC_I0(A_bar, A);
    not SMC_I1(B_bar, B);
    and SMC_I2(Z, A_bar, B_bar);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // NR2M6N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:11:39 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR2M8N(A, B, Z);
  input A, B;
  output Z;

    not SMC_I0(A_bar, A);
    not SMC_I1(B_bar, B);
    and SMC_I2(Z, A_bar, B_bar);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // NR2M8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:13:20 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module NR3B1M0N ( Z, B, C, NA );
   input B, C, NA;
   output Z;
      NR3B1M0N_UDP3(Z, B, C, NA);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc NA --> Z
    (NA => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // NR3B1M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:20:40 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module NR3B1M1N ( Z, B, C, NA );
   input B, C, NA;
   output Z;
      NR3B1M0N_UDP3(Z, B, C, NA);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc NA --> Z
    (NA => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // NR3B1M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:19:34 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module NR3B1M2N ( Z, B, C, NA );
   input B, C, NA;
   output Z;
      NR3B1M0N_UDP3(Z, B, C, NA);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc NA --> Z
    (NA => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // NR3B1M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:18:42 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module NR3B1M4N ( Z, B, C, NA );
   input B, C, NA;
   output Z;
      NR3B1M0N_UDP3(Z, B, C, NA);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc NA --> Z
    (NA => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // NR3B1M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:13:35 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module NR3M0N ( Z, A, B, C );
   input A, B, C;
   output Z;
      NR3M0N_UDP3(Z, A, B, C);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // NR3M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:14:10 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module NR3M1N ( Z, A, B, C );
   input A, B, C;
   output Z;
      NR3M0N_UDP3(Z, A, B, C);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // NR3M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:13:35 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module NR3M2N ( Z, A, B, C );
   input A, B, C;
   output Z;
      NR3M0N_UDP3(Z, A, B, C);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // NR3M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:11:54 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module NR3M4N ( Z, A, B, C );
   input A, B, C;
   output Z;
      NR3M0N_UDP3(Z, A, B, C);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // NR3M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:17:12 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module NR3M6N ( Z, A, B, C );
   input A, B, C;
   output Z;
      NR3M0N_UDP3(Z, A, B, C);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // NR3M6N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:16:16 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module NR3M8N ( Z, A, B, C );
   input A, B, C;
   output Z;
      NR3M0N_UDP3(Z, A, B, C);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // NR3M8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:16:03 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module NR4B1M0N ( Z, B, C, D, NA );
   input B, C, D, NA;
   output Z;
      NR4B1M0N_UDP4(Z, B, C, D, NA);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc D --> Z
    (D => Z) = (1.0, 1.0);

    // arc NA --> Z
    (NA => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // NR4B1M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:14:25 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module NR4B1M1N ( Z, B, C, D, NA );
   input B, C, D, NA;
   output Z;
      NR4B1M0N_UDP4(Z, B, C, D, NA);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc D --> Z
    (D => Z) = (1.0, 1.0);

    // arc NA --> Z
    (NA => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // NR4B1M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:13:50 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module NR4B1M2N ( Z, B, C, D, NA );
   input B, C, D, NA;
   output Z;
      NR4B1M0N_UDP4(Z, B, C, D, NA);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc D --> Z
    (D => Z) = (1.0, 1.0);

    // arc NA --> Z
    (NA => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // NR4B1M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:12:10 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module NR4B1M4N ( Z, B, C, D, NA );
   input B, C, D, NA;
   output Z;
      NR4B1M0N_UDP4(Z, B, C, D, NA);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc D --> Z
    (D => Z) = (1.0, 1.0);

    // arc NA --> Z
    (NA => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // NR4B1M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:17:27 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module NR4B2M0N ( Z, C, D, NA, NB );
   input C, D, NA, NB;
   output Z;
      NR4B2M0N_UDP4(Z, C, D, NA, NB);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc D --> Z
    (D => Z) = (1.0, 1.0);

    // arc NA --> Z
    (NA => Z) = (1.0, 1.0);

    // arc NB --> Z
    (NB => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // NR4B2M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:16:32 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module NR4B2M1N ( Z, C, D, NA, NB );
   input C, D, NA, NB;
   output Z;
      NR4B2M0N_UDP4(Z, C, D, NA, NB);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc D --> Z
    (D => Z) = (1.0, 1.0);

    // arc NA --> Z
    (NA => Z) = (1.0, 1.0);

    // arc NB --> Z
    (NB => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // NR4B2M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:13:50 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module NR4B2M2N ( Z, C, D, NA, NB );
   input C, D, NA, NB;
   output Z;
      NR4B2M0N_UDP4(Z, C, D, NA, NB);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc D --> Z
    (D => Z) = (1.0, 1.0);

    // arc NA --> Z
    (NA => Z) = (1.0, 1.0);

    // arc NB --> Z
    (NB => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // NR4B2M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:13:41 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module NR4B2M4N ( Z, C, D, NA, NB );
   input C, D, NA, NB;
   output Z;
      NR4B2M0N_UDP4(Z, C, D, NA, NB);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc D --> Z
    (D => Z) = (1.0, 1.0);

    // arc NA --> Z
    (NA => Z) = (1.0, 1.0);

    // arc NB --> Z
    (NB => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // NR4B2M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:14:40 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module NR4M0N ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;
      NR4M0N_UDP4(Z, A, B, C, D);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc D --> Z
    (D => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // NR4M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:13:42 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module NR4M1N ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;
      NR4M0N_UDP4(Z, A, B, C, D);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc D --> Z
    (D => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // NR4M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:12:24 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module NR4M2N ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;
      NR4M0N_UDP4(Z, A, B, C, D);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc D --> Z
    (D => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // NR4M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:14:05 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module NR4M4N ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;
      NR4M0N_UDP4(Z, A, B, C, D);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc D --> Z
    (D => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // NR4M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:14:40 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module NR4M6N ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;
      NR4M0N_UDP4(Z, A, B, C, D);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc D --> Z
    (D => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // NR4M6N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:17:12 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module NR4M8N ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;
      NR4M0N_UDP4(Z, A, B, C, D);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc D --> Z
    (D => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // NR4M8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:16:46 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA21M0N(A1, A2, B, Z);
  input A1, A2, B;
  output Z;

    and SMC_I0(OUT0, A1, B);
    and SMC_I1(OUT1, A2, B);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OA21M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:14:55 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA21M1N(A1, A2, B, Z);
  input A1, A2, B;
  output Z;

    and SMC_I0(OUT0, A1, B);
    and SMC_I1(OUT1, A2, B);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OA21M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:11:55 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA21M2N(A1, A2, B, Z);
  input A1, A2, B;
  output Z;

    and SMC_I0(OUT0, A1, B);
    and SMC_I1(OUT1, A2, B);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OA21M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:13:54 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA21M4N(A1, A2, B, Z);
  input A1, A2, B;
  output Z;

    and SMC_I0(OUT0, A1, B);
    and SMC_I1(OUT1, A2, B);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OA21M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:12:40 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA22M0N(A1, A2, B1, B2, Z);
  input A1, A2, B1, B2;
  output Z;

    and SMC_I0(OUT0, A2, B2);
    and SMC_I1(OUT1, A1, B2);
    and SMC_I2(OUT2, A1, B1);
    and SMC_I3(OUT3, A2, B1);
    or SMC_I4(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OA22M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:14:20 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA22M1N(A1, A2, B1, B2, Z);
  input A1, A2, B1, B2;
  output Z;

    and SMC_I0(OUT0, A2, B2);
    and SMC_I1(OUT1, A1, B2);
    and SMC_I2(OUT2, A1, B1);
    and SMC_I3(OUT3, A2, B1);
    or SMC_I4(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OA22M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:17:28 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA22M2N(A1, A2, B1, B2, Z);
  input A1, A2, B1, B2;
  output Z;

    and SMC_I0(OUT0, A2, B2);
    and SMC_I1(OUT1, A1, B2);
    and SMC_I2(OUT2, A1, B1);
    and SMC_I3(OUT3, A2, B1);
    or SMC_I4(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OA22M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:14:55 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA22M4N(A1, A2, B1, B2, Z);
  input A1, A2, B1, B2;
  output Z;

    and SMC_I0(OUT0, A2, B2);
    and SMC_I1(OUT1, A1, B2);
    and SMC_I2(OUT2, A1, B1);
    and SMC_I3(OUT3, A2, B1);
    or SMC_I4(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OA22M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:18:55 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI211B100M0N(A1, B, C, NA2, Z);
  input A1, B, C, NA2;
  output Z;

    not SMC_I0(C_bar, C);
    buf SMC_I1(OUT0, C_bar);
    not SMC_I2(B_bar, B);
    buf SMC_I3(OUT1, B_bar);
    not SMC_I4(A1_bar, A1);
    and SMC_I5(OUT2, A1_bar, NA2);
    or SMC_I6(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc NA2 --> Z
    (NA2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI211B100M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:20:01 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI211B100M1N(A1, B, C, NA2, Z);
  input A1, B, C, NA2;
  output Z;

    not SMC_I0(C_bar, C);
    buf SMC_I1(OUT0, C_bar);
    not SMC_I2(B_bar, B);
    buf SMC_I3(OUT1, B_bar);
    not SMC_I4(A1_bar, A1);
    and SMC_I5(OUT2, A1_bar, NA2);
    or SMC_I6(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc NA2 --> Z
    (NA2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI211B100M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:21:05 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI211B100M2N(A1, B, C, NA2, Z);
  input A1, B, C, NA2;
  output Z;

    not SMC_I0(C_bar, C);
    buf SMC_I1(OUT0, C_bar);
    not SMC_I2(B_bar, B);
    buf SMC_I3(OUT1, B_bar);
    not SMC_I4(A1_bar, A1);
    and SMC_I5(OUT2, A1_bar, NA2);
    or SMC_I6(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc NA2 --> Z
    (NA2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI211B100M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:14:41 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI211B100M4N(A1, B, C, NA2, Z);
  input A1, B, C, NA2;
  output Z;

    not SMC_I0(C_bar, C);
    buf SMC_I1(OUT0, C_bar);
    not SMC_I2(B_bar, B);
    buf SMC_I3(OUT1, B_bar);
    not SMC_I4(A1_bar, A1);
    and SMC_I5(OUT2, A1_bar, NA2);
    or SMC_I6(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc NA2 --> Z
    (NA2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI211B100M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:16:17 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI211M0N(A1, A2, B, C, Z);
  input A1, A2, B, C;
  output Z;

    not SMC_I0(C_bar, C);
    buf SMC_I1(OUT0, C_bar);
    not SMC_I2(A1_bar, A1);
    not SMC_I3(A2_bar, A2);
    and SMC_I4(OUT1, A1_bar, A2_bar);
    not SMC_I5(B_bar, B);
    buf SMC_I6(OUT2, B_bar);
    or SMC_I7(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI211M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:15:11 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI211M1N(A1, A2, B, C, Z);
  input A1, A2, B, C;
  output Z;

    not SMC_I0(C_bar, C);
    buf SMC_I1(OUT0, C_bar);
    not SMC_I2(A1_bar, A1);
    not SMC_I3(A2_bar, A2);
    and SMC_I4(OUT1, A1_bar, A2_bar);
    not SMC_I5(B_bar, B);
    buf SMC_I6(OUT2, B_bar);
    or SMC_I7(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI211M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:12:12 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI211M2N(A1, A2, B, C, Z);
  input A1, A2, B, C;
  output Z;

    not SMC_I0(C_bar, C);
    buf SMC_I1(OUT0, C_bar);
    not SMC_I2(A1_bar, A1);
    not SMC_I3(A2_bar, A2);
    and SMC_I4(OUT1, A1_bar, A2_bar);
    not SMC_I5(B_bar, B);
    buf SMC_I6(OUT2, B_bar);
    or SMC_I7(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI211M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:12:12 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI211M4N(A1, A2, B, C, Z);
  input A1, A2, B, C;
  output Z;

    not SMC_I0(C_bar, C);
    buf SMC_I1(OUT0, C_bar);
    not SMC_I2(A1_bar, A1);
    not SMC_I3(A2_bar, A2);
    and SMC_I4(OUT1, A1_bar, A2_bar);
    not SMC_I5(B_bar, B);
    buf SMC_I6(OUT2, B_bar);
    or SMC_I7(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI211M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:17:44 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21B01M0N(A1, A2, NB, Z);
  input A1, A2, NB;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(A2_bar, A2);
    and SMC_I2(OUT0, A1_bar, A2_bar);
    buf SMC_I3(OUT1, NB);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc NB --> Z
    (NB => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI21B01M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:15:12 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21B01M1N(A1, A2, NB, Z);
  input A1, A2, NB;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(A2_bar, A2);
    and SMC_I2(OUT0, A1_bar, A2_bar);
    buf SMC_I3(OUT1, NB);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc NB --> Z
    (NB => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI21B01M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:14:47 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21B01M2N(A1, A2, NB, Z);
  input A1, A2, NB;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(A2_bar, A2);
    and SMC_I2(OUT0, A1_bar, A2_bar);
    buf SMC_I3(OUT1, NB);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc NB --> Z
    (NB => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI21B01M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:14:37 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21B01M4N(A1, A2, NB, Z);
  input A1, A2, NB;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(A2_bar, A2);
    and SMC_I2(OUT0, A1_bar, A2_bar);
    buf SMC_I3(OUT1, NB);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc NB --> Z
    (NB => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI21B01M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:15:26 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21B10M0N(A1, B, NA2, Z);
  input A1, B, NA2;
  output Z;

    not SMC_I0(B_bar, B);
    buf SMC_I1(OUT0, B_bar);
    not SMC_I2(A1_bar, A1);
    and SMC_I3(OUT1, A1_bar, NA2);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc NA2 --> Z
    (NA2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI21B10M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:12:26 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21B10M1N(A1, B, NA2, Z);
  input A1, B, NA2;
  output Z;

    not SMC_I0(B_bar, B);
    buf SMC_I1(OUT0, B_bar);
    not SMC_I2(A1_bar, A1);
    and SMC_I3(OUT1, A1_bar, NA2);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc NA2 --> Z
    (NA2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI21B10M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:12:26 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21B10M2N(A1, B, NA2, Z);
  input A1, B, NA2;
  output Z;

    not SMC_I0(B_bar, B);
    buf SMC_I1(OUT0, B_bar);
    not SMC_I2(A1_bar, A1);
    and SMC_I3(OUT1, A1_bar, NA2);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc NA2 --> Z
    (NA2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI21B10M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:17:58 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21B10M4N(A1, B, NA2, Z);
  input A1, B, NA2;
  output Z;

    not SMC_I0(B_bar, B);
    buf SMC_I1(OUT0, B_bar);
    not SMC_I2(A1_bar, A1);
    and SMC_I3(OUT1, A1_bar, NA2);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc NA2 --> Z
    (NA2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI21B10M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:15:26 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21B20M0N(B, NA1, NA2, Z);
  input B, NA1, NA2;
  output Z;

    not SMC_I0(B_bar, B);
    buf SMC_I1(OUT0, B_bar);
    and SMC_I2(OUT1, NA1, NA2);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc NA1 --> Z
    (NA1 => Z) = (1.0, 1.0);

    // arc NA2 --> Z
    (NA2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI21B20M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:14:51 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21B20M1N(B, NA1, NA2, Z);
  input B, NA1, NA2;
  output Z;

    not SMC_I0(B_bar, B);
    buf SMC_I1(OUT0, B_bar);
    and SMC_I2(OUT1, NA1, NA2);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc NA1 --> Z
    (NA1 => Z) = (1.0, 1.0);

    // arc NA2 --> Z
    (NA2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI21B20M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:15:42 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21B20M2N(B, NA1, NA2, Z);
  input B, NA1, NA2;
  output Z;

    not SMC_I0(B_bar, B);
    buf SMC_I1(OUT0, B_bar);
    and SMC_I2(OUT1, NA1, NA2);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc NA1 --> Z
    (NA1 => Z) = (1.0, 1.0);

    // arc NA2 --> Z
    (NA2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI21B20M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:12:42 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21B20M4N(B, NA1, NA2, Z);
  input B, NA1, NA2;
  output Z;

    not SMC_I0(B_bar, B);
    buf SMC_I1(OUT0, B_bar);
    and SMC_I2(OUT1, NA1, NA2);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc NA1 --> Z
    (NA1 => Z) = (1.0, 1.0);

    // arc NA2 --> Z
    (NA2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI21B20M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:18:14 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21M0N(A1, A2, B, Z);
  input A1, A2, B;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(A2_bar, A2);
    and SMC_I2(OUT0, A1_bar, A2_bar);
    not SMC_I3(B_bar, B);
    buf SMC_I4(OUT1, B_bar);
    or SMC_I5(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI21M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:14:03 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21M1N(A1, A2, B, Z);
  input A1, A2, B;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(A2_bar, A2);
    and SMC_I2(OUT0, A1_bar, A2_bar);
    not SMC_I3(B_bar, B);
    buf SMC_I4(OUT1, B_bar);
    or SMC_I5(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI21M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:15:42 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21M2N(A1, A2, B, Z);
  input A1, A2, B;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(A2_bar, A2);
    and SMC_I2(OUT0, A1_bar, A2_bar);
    not SMC_I3(B_bar, B);
    buf SMC_I4(OUT1, B_bar);
    or SMC_I5(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI21M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:17:48 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21M3N(A1, A2, B, Z);
  input A1, A2, B;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(A2_bar, A2);
    and SMC_I2(OUT0, A1_bar, A2_bar);
    not SMC_I3(B_bar, B);
    buf SMC_I4(OUT1, B_bar);
    or SMC_I5(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI21M3N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:15:07 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21M4N(A1, A2, B, Z);
  input A1, A2, B;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(A2_bar, A2);
    and SMC_I2(OUT0, A1_bar, A2_bar);
    not SMC_I3(B_bar, B);
    buf SMC_I4(OUT1, B_bar);
    or SMC_I5(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI21M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:15:57 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21M6N(A1, A2, B, Z);
  input A1, A2, B;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(A2_bar, A2);
    and SMC_I2(OUT0, A1_bar, A2_bar);
    not SMC_I3(B_bar, B);
    buf SMC_I4(OUT1, B_bar);
    or SMC_I5(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI21M6N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:12:58 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21M8N(A1, A2, B, Z);
  input A1, A2, B;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(A2_bar, A2);
    and SMC_I2(OUT0, A1_bar, A2_bar);
    not SMC_I3(B_bar, B);
    buf SMC_I4(OUT1, B_bar);
    or SMC_I5(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI21M8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:15:58 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI221M0N ( Z, A1, A2, B1, B2, C );
   input A1, A2, B1, B2, C;
   output Z;
      OAI221M0N_UDP5(Z, A1, A2, B1, B2, C);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI221M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:17:37 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI221M1N ( Z, A1, A2, B1, B2, C );
   input A1, A2, B1, B2, C;
   output Z;
      OAI221M0N_UDP5(Z, A1, A2, B1, B2, C);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI221M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:18:30 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI221M2N ( Z, A1, A2, B1, B2, C );
   input A1, A2, B1, B2, C;
   output Z;
      OAI221M0N_UDP5(Z, A1, A2, B1, B2, C);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI221M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:16:14 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI221M4N ( Z, A1, A2, B1, B2, C );
   input A1, A2, B1, B2, C;
   output Z;
      OAI221M0N_UDP5(Z, A1, A2, B1, B2, C);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI221M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:17:53 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI222M0N ( Z, A1, A2, B1, B2, C1, C2 );
   input A1, A2, B1, B2, C1, C2;
   output Z;
      OAI222M0N_UDP6(Z, A1, A2, B1, B2, C1, C2);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);

    // arc C1 --> Z
    (C1 => Z) = (1.0, 1.0);

    // arc C2 --> Z
    (C2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI222M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:18:46 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI222M1N ( Z, A1, A2, B1, B2, C1, C2 );
   input A1, A2, B1, B2, C1, C2;
   output Z;
      OAI222M0N_UDP6(Z, A1, A2, B1, B2, C1, C2);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);

    // arc C1 --> Z
    (C1 => Z) = (1.0, 1.0);

    // arc C2 --> Z
    (C2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI222M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:16:14 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI222M2N ( Z, A1, A2, B1, B2, C1, C2 );
   input A1, A2, B1, B2, C1, C2;
   output Z;
      OAI222M0N_UDP6(Z, A1, A2, B1, B2, C1, C2);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);

    // arc C1 --> Z
    (C1 => Z) = (1.0, 1.0);

    // arc C2 --> Z
    (C2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI222M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:14:06 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI222M4N ( Z, A1, A2, B1, B2, C1, C2 );
   input A1, A2, B1, B2, C1, C2;
   output Z;
      OAI222M0N_UDP6(Z, A1, A2, B1, B2, C1, C2);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);

    // arc C1 --> Z
    (C1 => Z) = (1.0, 1.0);

    // arc C2 --> Z
    (C2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI222M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:17:53 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI22B10M0N ( Z, A1, B1, B2, NA2 );
   input A1, B1, B2, NA2;
   output Z;
      OAI22B10M0N_UDP4(Z, A1, B1, B2, NA2);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);

    // arc NA2 --> Z
    (NA2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI22B10M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:18:46 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI22B10M1N ( Z, A1, B1, B2, NA2 );
   input A1, B1, B2, NA2;
   output Z;
      OAI22B10M0N_UDP4(Z, A1, B1, B2, NA2);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);

    // arc NA2 --> Z
    (NA2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI22B10M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:14:05 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI22B10M2N ( Z, A1, B1, B2, NA2 );
   input A1, B1, B2, NA2;
   output Z;
      OAI22B10M0N_UDP4(Z, A1, B1, B2, NA2);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);

    // arc NA2 --> Z
    (NA2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI22B10M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:20:06 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI22B10M4N ( Z, A1, B1, B2, NA2 );
   input A1, B1, B2, NA2;
   output Z;
      OAI22B10M0N_UDP4(Z, A1, B1, B2, NA2);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);

    // arc NA2 --> Z
    (NA2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI22B10M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:16:28 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI22B20M0N ( Z, B1, B2, NA1, NA2 );
   input B1, B2, NA1, NA2;
   output Z;
      OAI22B20M0N_UDP4(Z, B1, B2, NA1, NA2);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);

    // arc NA1 --> Z
    (NA1 => Z) = (1.0, 1.0);

    // arc NA2 --> Z
    (NA2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI22B20M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:14:15 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI22B20M1N ( Z, B1, B2, NA1, NA2 );
   input B1, B2, NA1, NA2;
   output Z;
      OAI22B20M0N_UDP4(Z, B1, B2, NA1, NA2);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);

    // arc NA1 --> Z
    (NA1 => Z) = (1.0, 1.0);

    // arc NA2 --> Z
    (NA2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI22B20M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:18:07 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI22B20M2N ( Z, B1, B2, NA1, NA2 );
   input B1, B2, NA1, NA2;
   output Z;
      OAI22B20M0N_UDP4(Z, B1, B2, NA1, NA2);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);

    // arc NA1 --> Z
    (NA1 => Z) = (1.0, 1.0);

    // arc NA2 --> Z
    (NA2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI22B20M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:18:34 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI22B20M4N ( Z, B1, B2, NA1, NA2 );
   input B1, B2, NA1, NA2;
   output Z;
      OAI22B20M0N_UDP4(Z, B1, B2, NA1, NA2);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);

    // arc NA1 --> Z
    (NA1 => Z) = (1.0, 1.0);

    // arc NA2 --> Z
    (NA2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI22B20M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:16:37 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI22M0N ( Z, A1, A2, B1, B2 );
   input A1, A2, B1, B2;
   output Z;
      OAI22M0N_UDP4(Z, A1, A2, B1, B2);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI22M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:19:52 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI22M1N ( Z, A1, A2, B1, B2 );
   input A1, A2, B1, B2;
   output Z;
      OAI22M0N_UDP4(Z, A1, A2, B1, B2);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI22M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:15:10 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI22M2N ( Z, A1, A2, B1, B2 );
   input A1, A2, B1, B2;
   output Z;
      OAI22M0N_UDP4(Z, A1, A2, B1, B2);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI22M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:21:34 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI22M4N ( Z, A1, A2, B1, B2 );
   input A1, A2, B1, B2;
   output Z;
      OAI22M0N_UDP4(Z, A1, A2, B1, B2);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI22M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:17:23 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI31M0N ( Z, A1, A2, A3, B );
   input A1, A2, A3, B;
   output Z;
      OAI31M0N_UDP4(Z, A1, A2, A3, B);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc A3 --> Z
    (A3 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI31M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:18:24 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI31M1N ( Z, A1, A2, A3, B );
   input A1, A2, A3, B;
   output Z;
      OAI31M0N_UDP4(Z, A1, A2, A3, B);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc A3 --> Z
    (A3 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI31M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:18:52 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI31M2N ( Z, A1, A2, A3, B );
   input A1, A2, A3, B;
   output Z;
      OAI31M0N_UDP4(Z, A1, A2, A3, B);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc A3 --> Z
    (A3 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI31M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:19:10 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI31M4N ( Z, A1, A2, A3, B );
   input A1, A2, A3, B;
   output Z;
      OAI31M0N_UDP4(Z, A1, A2, A3, B);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc A3 --> Z
    (A3 => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI31M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:16:46 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI32M0N ( Z, A1, A2, A3, B1, B2 );
   input A1, A2, A3, B1, B2;
   output Z;
      OAI32M0N_UDP5(Z, A1, A2, A3, B1, B2);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc A3 --> Z
    (A3 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI32M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:19:18 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI32M1N ( Z, A1, A2, A3, B1, B2 );
   input A1, A2, A3, B1, B2;
   output Z;
      OAI32M0N_UDP5(Z, A1, A2, A3, B1, B2);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc A3 --> Z
    (A3 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI32M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:19:47 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI32M2N ( Z, A1, A2, A3, B1, B2 );
   input A1, A2, A3, B1, B2;
   output Z;
      OAI32M0N_UDP5(Z, A1, A2, A3, B1, B2);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc A3 --> Z
    (A3 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI32M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:20:51 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI32M4N ( Z, A1, A2, A3, B1, B2 );
   input A1, A2, A3, B1, B2;
   output Z;
      OAI32M0N_UDP5(Z, A1, A2, A3, B1, B2);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc A3 --> Z
    (A3 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI32M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:19:38 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI33M0N ( Z, A1, A2, A3, B1, B2, B3 );
   input A1, A2, A3, B1, B2, B3;
   output Z;
      OAI33M0N_UDP6(Z, A1, A2, A3, B1, B2, B3);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc A3 --> Z
    (A3 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);

    // arc B3 --> Z
    (B3 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI33M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:16:25 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI33M1N ( Z, A1, A2, A3, B1, B2, B3 );
   input A1, A2, A3, B1, B2, B3;
   output Z;
      OAI33M0N_UDP6(Z, A1, A2, A3, B1, B2, B3);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc A3 --> Z
    (A3 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);

    // arc B3 --> Z
    (B3 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI33M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:18:40 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI33M2N ( Z, A1, A2, A3, B1, B2, B3 );
   input A1, A2, A3, B1, B2, B3;
   output Z;
      OAI33M0N_UDP6(Z, A1, A2, A3, B1, B2, B3);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc A3 --> Z
    (A3 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);

    // arc B3 --> Z
    (B3 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI33M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:19:07 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI33M4N ( Z, A1, A2, A3, B1, B2, B3 );
   input A1, A2, A3, B1, B2, B3;
   output Z;
      OAI33M0N_UDP6(Z, A1, A2, A3, B1, B2, B3);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (1.0, 1.0);

    // arc A2 --> Z
    (A2 => Z) = (1.0, 1.0);

    // arc A3 --> Z
    (A3 => Z) = (1.0, 1.0);

    // arc B1 --> Z
    (B1 => Z) = (1.0, 1.0);

    // arc B2 --> Z
    (B2 => Z) = (1.0, 1.0);

    // arc B3 --> Z
    (B3 => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OAI33M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:19:33 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR2M0N(A, B, Z);
  input A, B;
  output Z;

    buf SMC_I0(OUT0, A);
    buf SMC_I1(OUT1, B);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OR2M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:17:01 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR2M1N(A, B, Z);
  input A, B;
  output Z;

    buf SMC_I0(OUT0, A);
    buf SMC_I1(OUT1, B);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OR2M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:20:03 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR2M2N(A, B, Z);
  input A, B;
  output Z;

    buf SMC_I0(OUT0, A);
    buf SMC_I1(OUT1, B);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OR2M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:21:39 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR2M4N(A, B, Z);
  input A, B;
  output Z;

    buf SMC_I0(OUT0, A);
    buf SMC_I1(OUT1, B);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OR2M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:14:02 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR2M6N(A, B, Z);
  input A, B;
  output Z;

    buf SMC_I0(OUT0, A);
    buf SMC_I1(OUT1, B);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OR2M6N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:14:03 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR2M8N(A, B, Z);
  input A, B;
  output Z;

    buf SMC_I0(OUT0, A);
    buf SMC_I1(OUT1, B);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OR2M8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:14:34 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR3M0N(A, B, C, Z);
  input A, B, C;
  output Z;

    buf SMC_I0(OUT0, B);
    buf SMC_I1(OUT1, A);
    buf SMC_I2(OUT2, C);
    or SMC_I3(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OR3M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:17:00 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR3M1N(A, B, C, Z);
  input A, B, C;
  output Z;

    buf SMC_I0(OUT0, B);
    buf SMC_I1(OUT1, A);
    buf SMC_I2(OUT2, C);
    or SMC_I3(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OR3M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:19:17 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR3M2N(A, B, C, Z);
  input A, B, C;
  output Z;

    buf SMC_I0(OUT0, B);
    buf SMC_I1(OUT1, A);
    buf SMC_I2(OUT2, C);
    or SMC_I3(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OR3M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:19:10 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR3M4N(A, B, C, Z);
  input A, B, C;
  output Z;

    buf SMC_I0(OUT0, B);
    buf SMC_I1(OUT1, A);
    buf SMC_I2(OUT2, C);
    or SMC_I3(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OR3M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:20:12 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR3M6N(A, B, C, Z);
  input A, B, C;
  output Z;

    buf SMC_I0(OUT0, B);
    buf SMC_I1(OUT1, A);
    buf SMC_I2(OUT2, C);
    or SMC_I3(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OR3M6N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:17:04 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR3M8N(A, B, C, Z);
  input A, B, C;
  output Z;

    buf SMC_I0(OUT0, B);
    buf SMC_I1(OUT1, A);
    buf SMC_I2(OUT2, C);
    or SMC_I3(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OR3M8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:20:16 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR4M0N(A, B, C, D, Z);
  input A, B, C, D;
  output Z;

    buf SMC_I0(OUT0, D);
    buf SMC_I1(OUT1, B);
    buf SMC_I2(OUT2, C);
    buf SMC_I3(OUT3, A);
    or SMC_I4(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc D --> Z
    (D => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OR4M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:14:14 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR4M1N(A, B, C, D, Z);
  input A, B, C, D;
  output Z;

    buf SMC_I0(OUT0, D);
    buf SMC_I1(OUT1, B);
    buf SMC_I2(OUT2, C);
    buf SMC_I3(OUT3, A);
    or SMC_I4(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc D --> Z
    (D => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OR4M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:20:43 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR4M2N(A, B, C, D, Z);
  input A, B, C, D;
  output Z;

    buf SMC_I0(OUT0, D);
    buf SMC_I1(OUT1, B);
    buf SMC_I2(OUT2, C);
    buf SMC_I3(OUT3, A);
    or SMC_I4(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc D --> Z
    (D => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OR4M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:14:59 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR4M4N(A, B, C, D, Z);
  input A, B, C, D;
  output Z;

    buf SMC_I0(OUT0, D);
    buf SMC_I1(OUT1, B);
    buf SMC_I2(OUT2, C);
    buf SMC_I3(OUT3, A);
    or SMC_I4(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc D --> Z
    (D => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OR4M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:17:44 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR4M6N(A, B, C, D, Z);
  input A, B, C, D;
  output Z;

    buf SMC_I0(OUT0, D);
    buf SMC_I1(OUT1, B);
    buf SMC_I2(OUT2, C);
    buf SMC_I3(OUT3, A);
    or SMC_I4(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc D --> Z
    (D => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OR4M6N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:14:48 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR4M8N(A, B, C, D, Z);
  input A, B, C, D;
  output Z;

    buf SMC_I0(OUT0, D);
    buf SMC_I1(OUT1, B);
    buf SMC_I2(OUT2, C);
    buf SMC_I3(OUT3, A);
    or SMC_I4(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc B --> Z
    (B => Z) = (1.0, 1.0);

    // arc C --> Z
    (C => Z) = (1.0, 1.0);

    // arc D --> Z
    (D => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // OR4M8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:21:52 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module REG1M1N(RD, RG, RGB, WE, RQB);
  input RD, RG, RGB, WE;
  output RQB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(RD), .en(WE), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(RD), .en(WE), .clear(1'b1), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(SMC_DINRQB, SMC_IQN);

    not SMC_I4(RGB_bar, RGB);
    nand SMC_I5(SMC_ZENRQB, RG, RGB_bar);


    bufif0 SMC_I6(RQB, SMC_DINRQB, SMC_ZENRQB);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc RD --> RQB
    (RD => RQB) = (1.0, 1.0);

    // arc RG --> RQB
    (RG => RQB) = (1.0,
        1.0,
        1.0,
        1.0,
        1.0,
        1.0);

    // arc RGB --> RQB
    (RGB => RQB) = (1.0,
        1.0,
        1.0,
        1.0,
        1.0,
        1.0);
        
    // arc RG --> RQB
    if (RD===1'b0 && WE===1'b0) 
        (RG => RQB) = (1.0, 1.0);
    if (RD===1'b1 && WE===1'b0) 
        (RG => RQB) = (1.0, 1.0);
    if (RD===1'b1 && WE===1'b1) 
        (RG => RQB) = (1.0, 1.0);

    // arc RGB --> RQB
    if (RD===1'b0 && WE===1'b0) 
        (RGB => RQB) = (1.0, 1.0);
    if (RD===1'b1 && WE===1'b0) 
        (RGB => RQB) = (1.0, 1.0);
    if (RD===1'b0 && WE===1'b1) 
        (RGB => RQB) = (1.0, 1.0);

    // arc WE --> RQB
    (posedge WE => ( RQB +: RD )) = (1.0, 1.0);
    
    // arc RG --> RQB
    if (WE===1'b1) 
        (RG => RQB) = (1.0, 1.0);

    // arc RGB --> RQB
    if (WE===1'b1) 
        (RGB => RQB) = (1.0, 1.0);
    
    // setup
    $setup( negedge RD, negedge WE , 1.0, notifier );

    // setup
    $setup( posedge RD, negedge WE , 1.0, notifier );

    // hold
    $hold( negedge WE, negedge RD, 1.0, notifier );

    // hold
    $hold( negedge WE, posedge RD, 1.0, notifier );

    // mpw
    $width( posedge WE, 1.0, 0, notifier );

    // mpw
    $width( negedge WE, 1.0, 0, notifier );

    $period( posedge WE, 0, notifier );
    $period( negedge WE, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // REG1M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:20:53 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module REG2M1N(RD, RG1, RG2, WE, RQ1B, RQ2B);
  input RD, RG1, RG2, WE;
  output RQ1B, RQ2B;
  reg notifier;

  wire SMC_LD_IN;
    not SMC_I0(SMC_LD_IN, RD);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(SMC_LD_IN), .en(WE), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(SMC_LD_IN), .en(WE), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(SMC_DINRQ1B, SMC_IQ);

    not SMC_I5(SMC_ZENRQ1B, RG1);


    bufif0 SMC_I6(RQ1B, SMC_DINRQ1B, SMC_ZENRQ1B);

    buf SMC_I7(SMC_DINRQ2B, SMC_IQ);

    not SMC_I8(SMC_ZENRQ2B, RG2);


    bufif0 SMC_I9(RQ2B, SMC_DINRQ2B, SMC_ZENRQ2B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc RD --> RQ1B
    (RD => RQ1B) = (1.0, 1.0);

    // arc RD --> RQ2B
    (RD => RQ2B) = (1.0, 1.0);

    // arc RG1 --> RQ1B
    (RG1 => RQ1B) = (1.0,
        1.0,
        1.0,
        1.0,
        1.0,
        1.0);

    // arc RG2 --> RQ2B
    (RG2 => RQ2B) = (1.0,
        1.0,
        1.0,
        1.0,
        1.0,
        1.0);

    // arc WE --> RQ1B
    (posedge WE => ( RQ1B -: RD )) = (1.0, 1.0);

    // arc WE --> RQ2B
    (posedge WE => ( RQ2B -: RD )) = (1.0, 1.0);



    // setup RD-hl WE-hl ()
    $setup(negedge RD, negedge WE, 1.0, notifier);

    // setup RD-lh WE-hl ()
    $setup(posedge RD, negedge WE, 1.0, notifier);

    // hold RD-hl WE-hl ()
    $hold(negedge WE, negedge RD, 1.0, notifier);

    // hold RD-lh WE-hl ()
    $hold(negedge WE, posedge RD, 1.0, notifier);

    // mpw WE-hl NS-hl ()
    $width(negedge WE, 1.0, 0, notifier);

    // mpw WE-lh NS-lh ()
    $width(posedge WE, 1.0, 0, notifier);

    $period( posedge WE, 0, notifier );
    $period( negedge WE, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // REG2M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:15:37 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module REGKM1N(RD, RQB);
  input RD;
  output RQB;

    buf(weak0,weak1) SMC_IO(RD, io_wire);
    buf              SMC_I1(io_wire, RD);
    not              SMC_I0(RQB, RD);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc RD --> RQB
    (RD => RQB) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // REGKM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:20:25 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module REGKM2N(RD, RQB);
  input RD;
  output RQB;

    not SMC_I0(RQB, RD);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc RD --> RQB
    (RD => RQB) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // REGKM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:15:08 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module REGKM4N(RD, RQB);
  input RD;
  output RQB;

    not SMC_I0(RQB, RD);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc RD --> RQB
    (RD => RQB) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // REGKM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:20:00 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFEM0N(D, E, SD, SE, CK, Q, QB);
  input D, E, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    SDFEM0N_UDP__OUT__ SMC_I1(SMC_NS_IN, D, E, SMC_IQ, SD, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(SE_bar, SE);
    and SMC_I7(shcheckCKDlh, E, SE_bar);

    not SMC_I8(shcheckCKElh, SE);

    buf SMC_I9(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup E-lh CK-lh (!SE)
    $setup(posedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // setup E-hl CK-lh (!SE)
    $setup(negedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (E&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (E&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold E-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        posedge E &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // hold E-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        negedge E &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (E&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (E&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFEM0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:15:04 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFEM1N(D, E, SD, SE, CK, Q, QB);
  input D, E, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    SDFEM0N_UDP__OUT__ SMC_I1(SMC_NS_IN, D, E, SMC_IQ, SD, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(SE_bar, SE);
    and SMC_I7(shcheckCKDlh, E, SE_bar);

    not SMC_I8(shcheckCKElh, SE);

    buf SMC_I9(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup E-lh CK-lh (!SE)
    $setup(posedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // setup E-hl CK-lh (!SE)
    $setup(negedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (E&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (E&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold E-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        posedge E &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // hold E-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        negedge E &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (E&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (E&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFEM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:17:56 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFEM2N(D, E, SD, SE, CK, Q, QB);
  input D, E, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    SDFEM0N_UDP__OUT__ SMC_I1(SMC_NS_IN, D, E, SMC_IQ, SD, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(SE_bar, SE);
    and SMC_I7(shcheckCKDlh, E, SE_bar);

    not SMC_I8(shcheckCKElh, SE);

    buf SMC_I9(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup E-lh CK-lh (!SE)
    $setup(posedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // setup E-hl CK-lh (!SE)
    $setup(negedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (E&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (E&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold E-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        posedge E &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // hold E-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        negedge E &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (E&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (E&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFEM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:22:06 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFEM4N(D, E, SD, SE, CK, Q, QB);
  input D, E, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    SDFEM0N_UDP__OUT__ SMC_I1(SMC_NS_IN, D, E, SMC_IQ, SD, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(SE_bar, SE);
    and SMC_I7(shcheckCKDlh, E, SE_bar);

    not SMC_I8(shcheckCKElh, SE);

    buf SMC_I9(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup E-lh CK-lh (!SE)
    $setup(posedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // setup E-hl CK-lh (!SE)
    $setup(negedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (E&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (E&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold E-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        posedge E &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // hold E-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        negedge E &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (E&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (E&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFEM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:16:54 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFEQBM0N(D, E, SD, SE, CK, QB);
  input D, E, SD, SE, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    SDFEQBM0N_UDP__OUT__ SMC_I1(SMC_NS_IN, D, E, SMC_IQ, SD, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(SE_bar, SE);
    and SMC_I6(shcheckCKDlh, E, SE_bar);

    not SMC_I7(shcheckCKElh, SE);

    buf SMC_I8(shcheckCKSDlh, SE);


  specify


    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup E-lh CK-lh (!SE)
    $setup(posedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // setup E-hl CK-lh (!SE)
    $setup(negedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (E&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (E&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold E-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        posedge E &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // hold E-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        negedge E &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (E&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (E&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFEQBM0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:14:30 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFEQBM1N(D, E, SD, SE, CK, QB);
  input D, E, SD, SE, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    SDFEQBM0N_UDP__OUT__ SMC_I1(SMC_NS_IN, D, E, SMC_IQ, SD, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(SE_bar, SE);
    and SMC_I6(shcheckCKDlh, E, SE_bar);

    not SMC_I7(shcheckCKElh, SE);

    buf SMC_I8(shcheckCKSDlh, SE);


  specify


    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup E-lh CK-lh (!SE)
    $setup(posedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // setup E-hl CK-lh (!SE)
    $setup(negedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (E&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (E&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold E-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        posedge E &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // hold E-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        negedge E &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (E&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (E&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFEQBM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:20:31 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFEQBM2N(D, E, SD, SE, CK, QB);
  input D, E, SD, SE, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    SDFEQBM0N_UDP__OUT__ SMC_I1(SMC_NS_IN, D, E, SMC_IQ, SD, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(SE_bar, SE);
    and SMC_I6(shcheckCKDlh, E, SE_bar);

    not SMC_I7(shcheckCKElh, SE);

    buf SMC_I8(shcheckCKSDlh, SE);


  specify


    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup E-lh CK-lh (!SE)
    $setup(posedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // setup E-hl CK-lh (!SE)
    $setup(negedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (E&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (E&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold E-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        posedge E &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // hold E-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        negedge E &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (E&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (E&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFEQBM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:15:14 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFEQBM4N(D, E, SD, SE, CK, QB);
  input D, E, SD, SE, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    SDFEQBM0N_UDP__OUT__ SMC_I1(SMC_NS_IN, D, E, SMC_IQ, SD, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(SE_bar, SE);
    and SMC_I6(shcheckCKDlh, E, SE_bar);

    not SMC_I7(shcheckCKElh, SE);

    buf SMC_I8(shcheckCKSDlh, SE);


  specify


    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup E-lh CK-lh (!SE)
    $setup(posedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // setup E-hl CK-lh (!SE)
    $setup(negedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (E&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (E&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold E-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        posedge E &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // hold E-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        negedge E &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (E&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (E&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFEQBM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:19:09 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFEZRM0N(D, E, RB, SD, SE, CK, Q, QB);
  input D, E, RB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    SDFEZRM0N_UDP__OUT__ SMC_I1(SMC_NS_IN, D, E, SMC_IQ, RB, SD, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(SE_bar, SE);
    and SMC_I7(shcheckCKDlh, E, RB, SE_bar);

    and SMC_I8(shcheckCKElh, RB, SE_bar);

    not SMC_I9(shcheckCKRBlh, SE);

    buf SMC_I10(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup E-hl CK-lh (RB&!SE)
    $setup(negedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // setup E-lh CK-lh (RB&!SE)
    $setup(posedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (E&RB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (E&RB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup RB-lh CK-lh (!SE)
    $setup(posedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // setup RB-hl CK-lh (!SE)
    $setup(negedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold E-hl CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        negedge E &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // hold E-lh CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        posedge E &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (E&RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (E&RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold RB-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        posedge RB &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // hold RB-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        negedge RB &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFEZRM0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:15:06 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFEZRM1N(D, E, RB, SD, SE, CK, Q, QB);
  input D, E, RB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    SDFEZRM0N_UDP__OUT__ SMC_I1(SMC_NS_IN, D, E, SMC_IQ, RB, SD, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(SE_bar, SE);
    and SMC_I7(shcheckCKDlh, E, RB, SE_bar);

    and SMC_I8(shcheckCKElh, RB, SE_bar);

    not SMC_I9(shcheckCKRBlh, SE);

    buf SMC_I10(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup E-hl CK-lh (RB&!SE)
    $setup(negedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // setup E-lh CK-lh (RB&!SE)
    $setup(posedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (E&RB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (E&RB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup RB-lh CK-lh (!SE)
    $setup(posedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // setup RB-hl CK-lh (!SE)
    $setup(negedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold E-hl CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        negedge E &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // hold E-lh CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        posedge E &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (E&RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (E&RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold RB-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        posedge RB &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // hold RB-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        negedge RB &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFEZRM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:20:02 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFEZRM2N(D, E, RB, SD, SE, CK, Q, QB);
  input D, E, RB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    SDFEZRM0N_UDP__OUT__ SMC_I1(SMC_NS_IN, D, E, SMC_IQ, RB, SD, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(SE_bar, SE);
    and SMC_I7(shcheckCKDlh, E, RB, SE_bar);

    and SMC_I8(shcheckCKElh, RB, SE_bar);

    not SMC_I9(shcheckCKRBlh, SE);

    buf SMC_I10(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup E-hl CK-lh (RB&!SE)
    $setup(negedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // setup E-lh CK-lh (RB&!SE)
    $setup(posedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (E&RB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (E&RB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup RB-lh CK-lh (!SE)
    $setup(posedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // setup RB-hl CK-lh (!SE)
    $setup(negedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold E-hl CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        negedge E &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // hold E-lh CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        posedge E &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (E&RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (E&RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold RB-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        posedge RB &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // hold RB-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        negedge RB &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFEZRM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:17:38 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFEZRM4N(D, E, RB, SD, SE, CK, Q, QB);
  input D, E, RB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    SDFEZRM0N_UDP__OUT__ SMC_I1(SMC_NS_IN, D, E, SMC_IQ, RB, SD, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(SE_bar, SE);
    and SMC_I7(shcheckCKDlh, E, RB, SE_bar);

    and SMC_I8(shcheckCKElh, RB, SE_bar);

    not SMC_I9(shcheckCKRBlh, SE);

    buf SMC_I10(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup E-hl CK-lh (RB&!SE)
    $setup(negedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // setup E-lh CK-lh (RB&!SE)
    $setup(posedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (E&RB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (E&RB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup RB-lh CK-lh (!SE)
    $setup(posedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // setup RB-hl CK-lh (!SE)
    $setup(negedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold E-hl CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        negedge E &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // hold E-lh CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        posedge E &&& (shcheckCKElh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (E&RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (E&RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold RB-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        posedge RB &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // hold RB-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        negedge RB &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFEZRM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:20:37 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFM0N(D, SD, SE, CK, Q, QB);
  input D, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(shcheckCKDlh, SE);

    buf SMC_I7(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFM0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:15:34 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFM1N(D, SD, SE, CK, Q, QB);
  input D, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(shcheckCKDlh, SE);

    buf SMC_I7(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:18:35 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFM2N(D, SD, SE, CK, Q, QB);
  input D, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(shcheckCKDlh, SE);

    buf SMC_I7(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:21:40 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFM4N(D, SD, SE, CK, Q, QB);
  input D, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(shcheckCKDlh, SE);

    buf SMC_I7(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:16:23 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQBM0N(D, SD, SE, CK, QB);
  input D, SD, SE, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(shcheckCKDlh, SE);

    buf SMC_I6(shcheckCKSDlh, SE);


  specify


    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQBM0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:20:20 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQBM1N(D, SD, SE, CK, QB);
  input D, SD, SE, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(shcheckCKDlh, SE);

    buf SMC_I6(shcheckCKSDlh, SE);


  specify


    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQBM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:21:17 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQBM2N(D, SD, SE, CK, QB);
  input D, SD, SE, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(shcheckCKDlh, SE);

    buf SMC_I6(shcheckCKSDlh, SE);


  specify


    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQBM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:18:07 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQBM4N(D, SD, SE, CK, QB);
  input D, SD, SE, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(shcheckCKDlh, SE);

    buf SMC_I6(shcheckCKSDlh, SE);


  specify


    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQBM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:21:49 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQBRM0N(D, RB, SD, SE, CK, QB);
  input D, RB, SD, SE, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(SE_bar, SE);
    and SMC_I6(shcheckCKDlh, RB, SE_bar);

    and SMC_I7(shcheckCKSDlh, RB, SE);

    buf SMC_I8(shcheckCKSElh, RB);


  specify


    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (RB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (RB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (RB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh (RB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (RB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (RB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 1.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQBRM0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:14:44 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQBRM1N(D, RB, SD, SE, CK, QB);
  input D, RB, SD, SE, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(SE_bar, SE);
    and SMC_I6(shcheckCKDlh, RB, SE_bar);

    and SMC_I7(shcheckCKSDlh, RB, SE);

    buf SMC_I8(shcheckCKSElh, RB);


  specify


    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (RB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (RB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (RB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh (RB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (RB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (RB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 1.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQBRM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:14:41 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQBRM2N(D, RB, SD, SE, CK, QB);
  input D, RB, SD, SE, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(SE_bar, SE);
    and SMC_I6(shcheckCKDlh, RB, SE_bar);

    and SMC_I7(shcheckCKSDlh, RB, SE);

    buf SMC_I8(shcheckCKSElh, RB);


  specify


    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (RB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (RB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (RB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh (RB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (RB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (RB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 1.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQBRM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:15:28 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQBRM4N(D, RB, SD, SE, CK, QB);
  input D, RB, SD, SE, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(SE_bar, SE);
    and SMC_I6(shcheckCKDlh, RB, SE_bar);

    and SMC_I7(shcheckCKSDlh, RB, SE);

    buf SMC_I8(shcheckCKSElh, RB);


  specify


    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (RB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (RB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (RB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh (RB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (RB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (RB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 1.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQBRM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:15:00 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQM0N(D, SD, SE, CK, Q);
  input D, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(shcheckCKDlh, SE);

    buf SMC_I5(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQM0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:22:05 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQM1N(D, SD, SE, CK, Q);
  input D, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(shcheckCKDlh, SE);

    buf SMC_I5(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:21:01 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQM2N(D, SD, SE, CK, Q);
  input D, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(shcheckCKDlh, SE);

    buf SMC_I5(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:15:44 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQM4N(D, SD, SE, CK, Q);
  input D, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(shcheckCKDlh, SE);

    buf SMC_I5(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:20:32 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQRM0N(D, RB, SD, SE, CK, Q);
  input D, RB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKDlh, RB, SE_bar);

    and SMC_I6(shcheckCKSDlh, RB, SE);

    buf SMC_I7(shcheckCKSElh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (RB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (RB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (RB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh (RB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (RB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (RB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 1.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQRM0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:19:39 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQRM1N(D, RB, SD, SE, CK, Q);
  input D, RB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKDlh, RB, SE_bar);

    and SMC_I6(shcheckCKSDlh, RB, SE);

    buf SMC_I7(shcheckCKSElh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (RB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (RB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (RB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh (RB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (RB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (RB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 1.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQRM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:22:50 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQRM2N(D, RB, SD, SE, CK, Q);
  input D, RB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKDlh, RB, SE_bar);

    and SMC_I6(shcheckCKSDlh, RB, SE);

    buf SMC_I7(shcheckCKSElh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (RB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (RB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (RB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh (RB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (RB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (RB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 1.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQRM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:21:49 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQRM4N(D, RB, SD, SE, CK, Q);
  input D, RB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKDlh, RB, SE_bar);

    and SMC_I6(shcheckCKSDlh, RB, SE);

    buf SMC_I7(shcheckCKSElh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (RB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (RB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (RB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh (RB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (RB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (RB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 1.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQRM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:18:20 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQSM0N(D, SB, SD, SE, CK, Q);
  input D, SB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(SB));

  `else // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(SB), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKDlh, SB, SE_bar);

    and SMC_I6(shcheckCKSDlh, SB, SE);

    buf SMC_I7(shcheckCKSElh, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (SB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (SB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (SB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh (SB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (SB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 1.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQSM0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:18:51 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQSM1N(D, SB, SD, SE, CK, Q);
  input D, SB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(SB));

  `else // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(SB), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKDlh, SB, SE_bar);

    and SMC_I6(shcheckCKSDlh, SB, SE);

    buf SMC_I7(shcheckCKSElh, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (SB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (SB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (SB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh (SB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (SB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 1.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQSM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:16:43 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQSM2N(D, SB, SD, SE, CK, Q);
  input D, SB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(SB));

  `else // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(SB), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKDlh, SB, SE_bar);

    and SMC_I6(shcheckCKSDlh, SB, SE);

    buf SMC_I7(shcheckCKSElh, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (SB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (SB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (SB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh (SB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (SB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 1.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQSM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:21:07 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQSM4N(D, SB, SD, SE, CK, Q);
  input D, SB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(SB));

  `else // functional //
    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(SB), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKDlh, SB, SE_bar);

    and SMC_I6(shcheckCKSDlh, SB, SE);

    buf SMC_I7(shcheckCKSElh, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (SB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (SB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (SB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh (SB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (SB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 1.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQSM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:16:02 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFRM0N(D, RB, SD, SE, CK, Q, QB);
  input D, RB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(SE_bar, SE);
    and SMC_I7(shcheckCKDlh, RB, SE_bar);

    and SMC_I8(shcheckCKSDlh, RB, SE);

    buf SMC_I9(shcheckCKSElh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (RB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (RB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (RB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh (RB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (RB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (RB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 1.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFRM0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:15:14 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFRM1N(D, RB, SD, SE, CK, Q, QB);
  input D, RB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(SE_bar, SE);
    and SMC_I7(shcheckCKDlh, RB, SE_bar);

    and SMC_I8(shcheckCKSDlh, RB, SE);

    buf SMC_I9(shcheckCKSElh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (RB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (RB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (RB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh (RB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (RB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (RB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 1.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFRM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:22:20 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFRM2N(D, RB, SD, SE, CK, Q, QB);
  input D, RB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(SE_bar, SE);
    and SMC_I7(shcheckCKDlh, RB, SE_bar);

    and SMC_I8(shcheckCKSDlh, RB, SE);

    buf SMC_I9(shcheckCKSElh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (RB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (RB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (RB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh (RB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (RB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (RB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 1.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFRM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:20:46 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFRM4N(D, RB, SD, SE, CK, Q, QB);
  input D, RB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(SE_bar, SE);
    and SMC_I7(shcheckCKDlh, RB, SE_bar);

    and SMC_I8(shcheckCKSDlh, RB, SE);

    buf SMC_I9(shcheckCKSElh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (RB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (RB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (RB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh (RB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (RB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (RB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 1.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFRM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:19:54 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFRSM0N(D, RB, SB, SD, SE, CK, Q, QB);
  input D, RB, SB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    inv_clr0 SMC_I0(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ));
  wire SMC_NS_IN;
    mux21 SMC_I2(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p1 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(SB));

  `else // functional //
    dff_p1 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I5(Q, SMC_IQ);

    buf SMC_I6(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I7(SE_bar, SE);
    and SMC_I8(shcheckCKDlh, RB, SB, SE_bar);

    buf SMC_I9(shcheckCKRBlh, SB);

    buf SMC_I10(shcheckCKSBlh, RB);

    and SMC_I11(shcheckCKSDlh, RB, SB, SE);

    and SMC_I12(shcheckCKSElh, RB, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (RB&SB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (RB&SB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SB-lh RB-lh ()
    $setup(posedge SB, posedge RB, 1.0, notifier);

    // setup SE-hl CK-lh (RB&SB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (RB&SB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (RB&SB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (RB&SB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB&SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB&SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SB-lh RB-lh ()
    $hold(posedge RB, posedge SB, 1.0, notifier);

    // hold SE-hl CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (RB&SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (RB&SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh (SB)
    $recovery(posedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh (RB)
    $recovery(posedge SB &&& (shcheckCKSBlh === 1'b1),
        posedge CK &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // removal RB-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        posedge RB &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // removal SB-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSBlh === 1'b1),
        posedge SB &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFRSM0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:21:16 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFRSM1N(D, RB, SB, SD, SE, CK, Q, QB);
  input D, RB, SB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    inv_clr0 SMC_I0(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ));
  wire SMC_NS_IN;
    mux21 SMC_I2(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p1 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(SB));

  `else // functional //
    dff_p1 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I5(Q, SMC_IQ);

    buf SMC_I6(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I7(SE_bar, SE);
    and SMC_I8(shcheckCKDlh, RB, SB, SE_bar);

    buf SMC_I9(shcheckCKRBlh, SB);

    buf SMC_I10(shcheckCKSBlh, RB);

    and SMC_I11(shcheckCKSDlh, RB, SB, SE);

    and SMC_I12(shcheckCKSElh, RB, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (RB&SB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (RB&SB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SB-lh RB-lh ()
    $setup(posedge SB, posedge RB, 1.0, notifier);

    // setup SE-hl CK-lh (RB&SB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (RB&SB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (RB&SB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (RB&SB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB&SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB&SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SB-lh RB-lh ()
    $hold(posedge RB, posedge SB, 1.0, notifier);

    // hold SE-hl CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (RB&SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (RB&SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh (SB)
    $recovery(posedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh (RB)
    $recovery(posedge SB &&& (shcheckCKSBlh === 1'b1),
        posedge CK &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // removal RB-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        posedge RB &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // removal SB-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSBlh === 1'b1),
        posedge SB &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFRSM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:15:16 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFRSM2N(D, RB, SB, SD, SE, CK, Q, QB);
  input D, RB, SB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    inv_clr0 SMC_I0(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ));
  wire SMC_NS_IN;
    mux21 SMC_I2(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p1 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(SB));

  `else // functional //
    dff_p1 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I5(Q, SMC_IQ);

    buf SMC_I6(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I7(SE_bar, SE);
    and SMC_I8(shcheckCKDlh, RB, SB, SE_bar);

    buf SMC_I9(shcheckCKRBlh, SB);

    buf SMC_I10(shcheckCKSBlh, RB);

    and SMC_I11(shcheckCKSDlh, RB, SB, SE);

    and SMC_I12(shcheckCKSElh, RB, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (RB&SB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (RB&SB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SB-lh RB-lh ()
    $setup(posedge SB, posedge RB, 1.0, notifier);

    // setup SE-hl CK-lh (RB&SB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (RB&SB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (RB&SB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (RB&SB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB&SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB&SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SB-lh RB-lh ()
    $hold(posedge RB, posedge SB, 1.0, notifier);

    // hold SE-hl CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (RB&SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (RB&SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh (SB)
    $recovery(posedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh (RB)
    $recovery(posedge SB &&& (shcheckCKSBlh === 1'b1),
        posedge CK &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // removal RB-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        posedge RB &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // removal SB-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSBlh === 1'b1),
        posedge SB &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFRSM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:23:13 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFRSM4N(D, RB, SB, SD, SE, CK, Q, QB);
  input D, RB, SB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    inv_clr0 SMC_I0(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ));
  wire SMC_NS_IN;
    mux21 SMC_I2(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p1 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
        .preset(SB));

  `else // functional //
    dff_p1 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB), .preset(SB),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I5(Q, SMC_IQ);

    buf SMC_I6(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I7(SE_bar, SE);
    and SMC_I8(shcheckCKDlh, RB, SB, SE_bar);

    buf SMC_I9(shcheckCKRBlh, SB);

    buf SMC_I10(shcheckCKSBlh, RB);

    and SMC_I11(shcheckCKSDlh, RB, SB, SE);

    and SMC_I12(shcheckCKSElh, RB, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (1.0, 1.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (RB&SB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (RB&SB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SB-lh RB-lh ()
    $setup(posedge SB, posedge RB, 1.0, notifier);

    // setup SE-hl CK-lh (RB&SB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (RB&SB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (RB&SB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (RB&SB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (RB&SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (RB&SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SB-lh RB-lh ()
    $hold(posedge RB, posedge SB, 1.0, notifier);

    // hold SE-hl CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (RB&SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (RB&SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (RB&SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery RB-lh CK-lh (SB)
    $recovery(posedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh (RB)
    $recovery(posedge SB &&& (shcheckCKSBlh === 1'b1),
        posedge CK &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // removal RB-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        posedge RB &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // removal SB-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSBlh === 1'b1),
        posedge SB &&& (shcheckCKSBlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFRSM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:17:00 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFSM0N(D, SB, SD, SE, CK, Q, QB);
  input D, SB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p1 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(SB));

  `else // functional //
    dff_p1 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(SB), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(SE_bar, SE);
    and SMC_I7(shcheckCKDlh, SB, SE_bar);

    and SMC_I8(shcheckCKSDlh, SB, SE);

    buf SMC_I9(shcheckCKSElh, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (SB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (SB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (SB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh (SB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (SB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 1.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFSM0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:19:23 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFSM1N(D, SB, SD, SE, CK, Q, QB);
  input D, SB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p1 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(SB));

  `else // functional //
    dff_p1 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(SB), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(SE_bar, SE);
    and SMC_I7(shcheckCKDlh, SB, SE_bar);

    and SMC_I8(shcheckCKSDlh, SB, SE);

    buf SMC_I9(shcheckCKSElh, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (SB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (SB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (SB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh (SB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (SB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 1.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFSM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:22:01 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFSM2N(D, SB, SD, SE, CK, Q, QB);
  input D, SB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p1 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(SB));

  `else // functional //
    dff_p1 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(SB), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(SE_bar, SE);
    and SMC_I7(shcheckCKDlh, SB, SE_bar);

    and SMC_I8(shcheckCKSDlh, SB, SE);

    buf SMC_I9(shcheckCKSElh, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (SB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (SB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (SB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh (SB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (SB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 1.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFSM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:21:09 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFSM4N(D, SB, SD, SE, CK, Q, QB);
  input D, SB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //
    dff_p1 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(SB));

  `else // functional //
    dff_p1 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(SB), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(SE_bar, SE);
    and SMC_I7(shcheckCKDlh, SB, SE_bar);

    and SMC_I8(shcheckCKSDlh, SB, SE);

    buf SMC_I9(shcheckCKSElh, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (1.0, 1.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl CK-lh (SB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-lh CK-lh (SB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup SE-lh CK-lh (SB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh (SB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // setup SD-hl CK-lh (SB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (SB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold SE-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 1.0, notifier);

    // hold SD-hl CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 1.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFSM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:21:43 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFZRM0N(D, RB, SD, SE, CK, Q, QB);
  input D, RB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    and SMC_I1(OUT0, SD, SE);
    not SMC_I2(SE_bar, SE);
    and SMC_I3(OUT1, D, RB, SE_bar);
    or SMC_I4(SMC_NS_IN, OUT0, OUT1);


  `ifdef functional // functional //
    dff_p0 SMC_I5(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I5(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I7(Q, SMC_IQ);

    buf SMC_I8(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I9(shcheckCKDlh, SE);

    not SMC_I10(shcheckCKRBlh, SE);

    buf SMC_I11(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup RB-hl CK-lh (!SE)
    $setup(negedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // setup RB-lh CK-lh (!SE)
    $setup(posedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold RB-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        negedge RB &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // hold RB-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        posedge RB &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFZRM0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:16:38 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFZRM1N(D, RB, SD, SE, CK, Q, QB);
  input D, RB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    and SMC_I1(OUT0, SD, SE);
    not SMC_I2(SE_bar, SE);
    and SMC_I3(OUT1, D, RB, SE_bar);
    or SMC_I4(SMC_NS_IN, OUT0, OUT1);


  `ifdef functional // functional //
    dff_p0 SMC_I5(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I5(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I7(Q, SMC_IQ);

    buf SMC_I8(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I9(shcheckCKDlh, SE);

    not SMC_I10(shcheckCKRBlh, SE);

    buf SMC_I11(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup RB-hl CK-lh (!SE)
    $setup(negedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // setup RB-lh CK-lh (!SE)
    $setup(posedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold RB-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        negedge RB &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // hold RB-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        posedge RB &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFZRM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:22:45 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFZRM2N(D, RB, SD, SE, CK, Q, QB);
  input D, RB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    and SMC_I1(OUT0, SD, SE);
    not SMC_I2(SE_bar, SE);
    and SMC_I3(OUT1, D, RB, SE_bar);
    or SMC_I4(SMC_NS_IN, OUT0, OUT1);


  `ifdef functional // functional //
    dff_p0 SMC_I5(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I5(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I7(Q, SMC_IQ);

    buf SMC_I8(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I9(shcheckCKDlh, SE);

    not SMC_I10(shcheckCKRBlh, SE);

    buf SMC_I11(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup RB-hl CK-lh (!SE)
    $setup(negedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // setup RB-lh CK-lh (!SE)
    $setup(posedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold RB-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        negedge RB &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // hold RB-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        posedge RB &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFZRM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:16:49 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFZRM4N(D, RB, SD, SE, CK, Q, QB);
  input D, RB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    and SMC_I1(OUT0, SD, SE);
    not SMC_I2(SE_bar, SE);
    and SMC_I3(OUT1, D, RB, SE_bar);
    or SMC_I4(SMC_NS_IN, OUT0, OUT1);


  `ifdef functional // functional //
    dff_p0 SMC_I5(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    dff_p0 SMC_I5(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I7(Q, SMC_IQ);

    buf SMC_I8(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I9(shcheckCKDlh, SE);

    not SMC_I10(shcheckCKRBlh, SE);

    buf SMC_I11(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (1.0, 1.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (1.0, 1.0);



    // setup D-lh CK-lh (!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup D-hl CK-lh (!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // setup RB-hl CK-lh (!SE)
    $setup(negedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // setup RB-lh CK-lh (!SE)
    $setup(posedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 1.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 1.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold D-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold D-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 1.0, notifier);

    // hold RB-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        negedge RB &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // hold RB-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        posedge RB &&& (shcheckCKRBlh === 1'b1), 1.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 1.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 1.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 1.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 1.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 1.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFZRM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:23:53 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module TIE0N(Z);
  output Z;

    buf SMC_I0(Z, 1'b0);


  `ifdef functional // functional //

  `else // functional //

  specify




  endspecify

  `endif // functional //
endmodule     // TIE0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:19:13 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module TIE1N(Z);
  output Z;

    buf SMC_I0(Z, 1'b1);


  `ifdef functional // functional //

  `else // functional //

  specify




  endspecify

  `endif // functional //
endmodule     // TIE1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:21:02 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module XNR2M0N(A, B, Z);
  input A, B;
  output Z;

    xnor SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
     if ( A===1'b1 )
    ( posedge A => ( Z +: A ) ) = (1.0, 1.0);
     if ( A===1'b0 )
    ( negedge A => ( Z +: A ) ) = (1.0, 1.0);

    // arc B --> Z
     if ( B===1'b1 )
    ( posedge B => ( Z +: B ) ) = (1.0, 1.0);
     if ( B===1'b0 )
    ( negedge B => ( Z +: B ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // XNR2M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:16:54 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module XNR2M1N(A, B, Z);
  input A, B;
  output Z;

    xnor SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
     if ( A===1'b1 )
    ( posedge A => ( Z +: A ) ) = (1.0, 1.0);
     if ( A===1'b0 )
    ( negedge A => ( Z +: A ) ) = (1.0, 1.0);

    // arc B --> Z
     if ( B===1'b1 )
    ( posedge B => ( Z +: B ) ) = (1.0, 1.0);
     if ( B===1'b0 )
    ( negedge B => ( Z +: B ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // XNR2M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:22:35 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module XNR2M2N(A, B, Z);
  input A, B;
  output Z;

    xnor SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
     if ( A===1'b1 )
    ( posedge A => ( Z +: A ) ) = (1.0, 1.0);
     if ( A===1'b0 )
    ( negedge A => ( Z +: A ) ) = (1.0, 1.0);

    // arc B --> Z
     if ( B===1'b1 )
    ( posedge B => ( Z +: B ) ) = (1.0, 1.0);
     if ( B===1'b0 )
    ( negedge B => ( Z +: B ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // XNR2M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:16:55 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module XNR2M4N(A, B, Z);
  input A, B;
  output Z;

    xnor SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
     if ( A===1'b1 )
    ( posedge A => ( Z +: A ) ) = (1.0, 1.0);
     if ( A===1'b0 )
    ( negedge A => ( Z +: A ) ) = (1.0, 1.0);

    // arc B --> Z
     if ( B===1'b1 )
    ( posedge B => ( Z +: B ) ) = (1.0, 1.0);
     if ( B===1'b0 )
    ( negedge B => ( Z +: B ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // XNR2M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:16:14 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module XNR3M0N ( Z, A, B, C );
   input A, B, C;
   output Z;
      XNR3M0N_UDP3(Z, A, B, C);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        ( posedge A => ( Z +: A ) ) = (1.0, 1.0);
        ( negedge A => ( Z +: A ) ) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        ( posedge B => ( Z +: B ) ) = (1.0, 1.0);
        ( negedge B => ( Z +: B ) ) = (1.0, 1.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1) 
        (C => Z) = (1.0, 1.0);
    ifnone
        ( posedge C => ( Z +: C ) ) = (1.0, 1.0);
        ( negedge C => ( Z +: C ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // XNR3M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:19:51 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module XNR3M1N ( Z, A, B, C );
   input A, B, C;
   output Z;
      XNR3M0N_UDP3(Z, A, B, C);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        ( posedge A => ( Z +: A ) ) = (1.0, 1.0);
        ( negedge A => ( Z +: A ) ) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        ( posedge B => ( Z +: B ) ) = (1.0, 1.0);
        ( negedge B => ( Z +: B ) ) = (1.0, 1.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1) 
        (C => Z) = (1.0, 1.0);
    ifnone
        ( posedge C => ( Z +: C ) ) = (1.0, 1.0);
        ( negedge C => ( Z +: C ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // XNR3M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:21:16 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module XNR3M2N ( Z, A, B, C );
   input A, B, C;
   output Z;
      XNR3M0N_UDP3(Z, A, B, C);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        ( posedge A => ( Z +: A ) ) = (1.0, 1.0);
        ( negedge A => ( Z +: A ) ) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        ( posedge B => ( Z +: B ) ) = (1.0, 1.0);
        ( negedge B => ( Z +: B ) ) = (1.0, 1.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1) 
        (C => Z) = (1.0, 1.0);
    ifnone
        ( posedge C => ( Z +: C ) ) = (1.0, 1.0);
        ( negedge C => ( Z +: C ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // XNR3M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:20:23 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module XNR3M4N ( Z, A, B, C );
   input A, B, C;
   output Z;
      XNR3M0N_UDP3(Z, A, B, C);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        ( posedge A => ( Z +: A ) ) = (1.0, 1.0);
        ( negedge A => ( Z +: A ) ) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        ( posedge B => ( Z +: B ) ) = (1.0, 1.0);
        ( negedge B => ( Z +: B ) ) = (1.0, 1.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1) 
        (C => Z) = (1.0, 1.0);
    ifnone
        ( posedge C => ( Z +: C ) ) = (1.0, 1.0);
        ( negedge C => ( Z +: C ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // XNR3M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 14:48:47 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module XOR2M0N(A, B, Z);
  input A, B;
  output Z;

    xor SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
     if ( A===1'b1 )
    ( posedge A => ( Z +: A ) ) = (1.0, 1.0);
     if ( A===1'b0 )
    ( negedge A => ( Z +: A ) ) = (1.0, 1.0);

    // arc B --> Z
     if ( B===1'b1 )
    ( posedge B => ( Z +: B ) ) = (1.0, 1.0);
     if ( B===1'b0 )
    ( negedge B => ( Z +: B ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // XOR2M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:20:50 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module XOR2M1N(A, B, Z);
  input A, B;
  output Z;

    xor SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
     if ( A===1'b1 )
    ( posedge A => ( Z +: A ) ) = (1.0, 1.0);
     if ( A===1'b0 )
    ( negedge A => ( Z +: A ) ) = (1.0, 1.0);

    // arc B --> Z
     if ( B===1'b1 )
    ( posedge B => ( Z +: B ) ) = (1.0, 1.0);
     if ( B===1'b0 )
    ( negedge B => ( Z +: B ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // XOR2M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:16:56 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module XOR2M2N(A, B, Z);
  input A, B;
  output Z;

    xor SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
     if ( A===1'b1 )
    ( posedge A => ( Z +: A ) ) = (1.0, 1.0);
     if ( A===1'b0 )
    ( negedge A => ( Z +: A ) ) = (1.0, 1.0);

    // arc B --> Z
     if ( B===1'b1 )
    ( posedge B => ( Z +: B ) ) = (1.0, 1.0);
     if ( B===1'b0 )
    ( negedge B => ( Z +: B ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // XOR2M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:16:57 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module XOR2M3N(A, B, Z);
  input A, B;
  output Z;

    xor SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
     if ( A===1'b1 )
    ( posedge A => ( Z +: A ) ) = (1.0, 1.0);
     if ( A===1'b0 )
    ( negedge A => ( Z +: A ) ) = (1.0, 1.0);

    // arc B --> Z
     if ( B===1'b1 )
    ( posedge B => ( Z +: B ) ) = (1.0, 1.0);
     if ( B===1'b0 )
    ( negedge B => ( Z +: B ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // XOR2M3N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:21:46 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module XOR2M4N(A, B, Z);
  input A, B;
  output Z;

    xor SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
     if ( A===1'b1 )
    ( posedge A => ( Z +: A ) ) = (1.0, 1.0);
     if ( A===1'b0 )
    ( negedge A => ( Z +: A ) ) = (1.0, 1.0);

    // arc B --> Z
     if ( B===1'b1 )
    ( posedge B => ( Z +: B ) ) = (1.0, 1.0);
     if ( B===1'b0 )
    ( negedge B => ( Z +: B ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // XOR2M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:16:29 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module XOR2M8N(A, B, Z);
  input A, B;
  output Z;

    xor SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
     if ( A===1'b1 )
    ( posedge A => ( Z +: A ) ) = (1.0, 1.0);
     if ( A===1'b0 )
    ( negedge A => ( Z +: A ) ) = (1.0, 1.0);

    // arc B --> Z
     if ( B===1'b1 )
    ( posedge B => ( Z +: B ) ) = (1.0, 1.0);
     if ( B===1'b0 )
    ( negedge B => ( Z +: B ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // XOR2M8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Mon Aug  1 19:11:58 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module XOR3M0N ( Z, A, B, C );
   input A, B, C;
   output Z;
      XOR3M0N_UDP3(Z, A, B, C);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        ( posedge A => ( Z +: A ) ) = (1.0, 1.0);
        ( negedge A => ( Z +: A ) ) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        ( posedge B => ( Z +: B ) ) = (1.0, 1.0);
        ( negedge B => ( Z +: B ) ) = (1.0, 1.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1) 
        (C => Z) = (1.0, 1.0);
    ifnone
        ( posedge C => ( Z +: C ) ) = (1.0, 1.0);
        ( negedge C => ( Z +: C ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // XOR3M0N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:22:00 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module XOR3M1N ( Z, A, B, C );
   input A, B, C;
   output Z;
      XOR3M0N_UDP3(Z, A, B, C);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        ( posedge A => ( Z +: A ) ) = (1.0, 1.0);
        ( negedge A => ( Z +: A ) ) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        ( posedge B => ( Z +: B ) ) = (1.0, 1.0);
        ( negedge B => ( Z +: B ) ) = (1.0, 1.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1) 
        (C => Z) = (1.0, 1.0);
    ifnone
        ( posedge C => ( Z +: C ) ) = (1.0, 1.0);
        ( negedge C => ( Z +: C ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // XOR3M1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:21:31 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module XOR3M2N ( Z, A, B, C );
   input A, B, C;
   output Z;
      XOR3M0N_UDP3(Z, A, B, C);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        ( posedge A => ( Z +: A ) ) = (1.0, 1.0);
        ( negedge A => ( Z +: A ) ) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        ( posedge B => ( Z +: B ) ) = (1.0, 1.0);
        ( negedge B => ( Z +: B ) ) = (1.0, 1.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1) 
        (C => Z) = (1.0, 1.0);
    ifnone
        ( posedge C => ( Z +: C ) ) = (1.0, 1.0);
        ( negedge C => ( Z +: C ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // XOR3M2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:20:38 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine 
module XOR3M4N ( Z, A, B, C );
   input A, B, C;
   output Z;
      XOR3M0N_UDP3(Z, A, B, C);
   
  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b0 && C===1'b1) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b0) 
        (A => Z) = (1.0, 1.0);
    if (B===1'b1 && C===1'b1) 
        (A => Z) = (1.0, 1.0);
    ifnone
        ( posedge A => ( Z +: A ) ) = (1.0, 1.0);
        ( negedge A => ( Z +: A ) ) = (1.0, 1.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b0 && C===1'b1) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b0) 
        (B => Z) = (1.0, 1.0);
    if (A===1'b1 && C===1'b1) 
        (B => Z) = (1.0, 1.0);
    ifnone
        ( posedge B => ( Z +: B ) ) = (1.0, 1.0);
        ( negedge B => ( Z +: B ) ) = (1.0, 1.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b0 && B===1'b1) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b0) 
        (C => Z) = (1.0, 1.0);
    if (A===1'b1 && B===1'b1) 
        (C => Z) = (1.0, 1.0);
    ifnone
        ( posedge C => ( Z +: C ) ) = (1.0, 1.0);
        ( negedge C => ( Z +: C ) ) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // XOR3M4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 21:11:24 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ISHM12N(A, E, Z);
  input A, E;
  output Z;

    buf SMC_I0(OUT0, A);
    buf SMC_I1(OUT1, E);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc E --> Z
    (E => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ISHM12N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 21:11:23 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ISHM16N(A, E, Z);
  input A, E;
  output Z;

    buf SMC_I0(OUT0, A);
    buf SMC_I1(OUT1, E);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc E --> Z
    (E => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ISHM16N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 21:16:58 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ISHM1N(A, E, Z);
  input A, E;
  output Z;

    buf SMC_I0(OUT0, A);
    buf SMC_I1(OUT1, E);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc E --> Z
    (E => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ISHM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 07:18:30 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ISHM20N(A, E, Z);
  input A, E;
  output Z;

    buf SMC_I0(OUT0, A);
    buf SMC_I1(OUT1, E);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc E --> Z
    (E => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ISHM20N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 07:13:52 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ISHM2N(A, E, Z);
  input A, E;
  output Z;

    buf SMC_I0(OUT0, A);
    buf SMC_I1(OUT1, E);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc E --> Z
    (E => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ISHM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 07:13:53 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ISHM32N(A, E, Z);
  input A, E;
  output Z;

    buf SMC_I0(OUT0, A);
    buf SMC_I1(OUT1, E);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc E --> Z
    (E => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ISHM32N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 21:16:59 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ISHM3N(A, E, Z);
  input A, E;
  output Z;

    buf SMC_I0(OUT0, A);
    buf SMC_I1(OUT1, E);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc E --> Z
    (E => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ISHM3N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 07:16:05 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ISHM4N(A, E, Z);
  input A, E;
  output Z;

    buf SMC_I0(OUT0, A);
    buf SMC_I1(OUT1, E);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc E --> Z
    (E => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ISHM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 21:11:20 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ISHM6N(A, E, Z);
  input A, E;
  output Z;

    buf SMC_I0(OUT0, A);
    buf SMC_I1(OUT1, E);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc E --> Z
    (E => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ISHM6N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 21:16:38 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ISHM8N(A, E, Z);
  input A, E;
  output Z;

    buf SMC_I0(OUT0, A);
    buf SMC_I1(OUT1, E);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc E --> Z
    (E => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ISHM8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 07:17:26 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ISLM12N(A, E, Z);
  input A, E;
  output Z;

    not SMC_I0(E_bar, E);
    and SMC_I1(Z, A, E_bar);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc E --> Z
    (E => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ISLM12N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 07:14:28 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ISLM16N(A, E, Z);
  input A, E;
  output Z;

    not SMC_I0(E_bar, E);
    and SMC_I1(Z, A, E_bar);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc E --> Z
    (E => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ISLM16N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 21:11:23 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ISLM1N(A, E, Z);
  input A, E;
  output Z;

    not SMC_I0(E_bar, E);
    and SMC_I1(Z, A, E_bar);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc E --> Z
    (E => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ISLM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 07:17:32 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ISLM20N(A, E, Z);
  input A, E;
  output Z;

    not SMC_I0(E_bar, E);
    and SMC_I1(Z, A, E_bar);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc E --> Z
    (E => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ISLM20N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 07:16:08 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ISLM2N(A, E, Z);
  input A, E;
  output Z;

    not SMC_I0(E_bar, E);
    and SMC_I1(Z, A, E_bar);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc E --> Z
    (E => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ISLM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 07:18:35 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ISLM32N(A, E, Z);
  input A, E;
  output Z;

    not SMC_I0(E_bar, E);
    and SMC_I1(Z, A, E_bar);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc E --> Z
    (E => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ISLM32N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 07:14:26 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ISLM3N(A, E, Z);
  input A, E;
  output Z;

    not SMC_I0(E_bar, E);
    and SMC_I1(Z, A, E_bar);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc E --> Z
    (E => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ISLM3N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 21:16:35 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ISLM4N(A, E, Z);
  input A, E;
  output Z;

    not SMC_I0(E_bar, E);
    and SMC_I1(Z, A, E_bar);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc E --> Z
    (E => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ISLM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 07:14:27 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ISLM6N(A, E, Z);
  input A, E;
  output Z;

    not SMC_I0(E_bar, E);
    and SMC_I1(Z, A, E_bar);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc E --> Z
    (E => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ISLM6N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 21:11:23 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ISLM8N(A, E, Z);
  input A, E;
  output Z;

    not SMC_I0(E_bar, E);
    and SMC_I1(Z, A, E_bar);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);

    // arc E --> Z
    (E => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // ISLM8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 07:17:29 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LALM12N(D, G, Q, QB);
  input D, G;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc D --> Q
    (D => Q) = (1.0, 1.0);

    // arc D --> QB
    (D => QB) = (1.0, 1.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (1.0, 1.0);

    // arc G --> QB
    (posedge G => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl G-hl ()
    $setup(negedge D, negedge G, 1.0, notifier);

    // setup D-lh G-hl ()
    $setup(posedge D, negedge G, 1.0, notifier);

    // hold D-hl G-hl ()
    $hold(negedge G, negedge D, 1.0, notifier);

    // hold D-lh G-hl ()
    $hold(negedge G, posedge D, 1.0, notifier);

    // mpw G-hl NS-hl ()
    $width(negedge G, 1.0, 0, notifier);

    // mpw G-lh NS-lh ()
    $width(posedge G, 1.0, 0, notifier);

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LALM12N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 21:11:30 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LALM16N(D, G, Q, QB);
  input D, G;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc D --> Q
    (D => Q) = (1.0, 1.0);

    // arc D --> QB
    (D => QB) = (1.0, 1.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (1.0, 1.0);

    // arc G --> QB
    (posedge G => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl G-hl ()
    $setup(negedge D, negedge G, 1.0, notifier);

    // setup D-lh G-hl ()
    $setup(posedge D, negedge G, 1.0, notifier);

    // hold D-hl G-hl ()
    $hold(negedge G, negedge D, 1.0, notifier);

    // hold D-lh G-hl ()
    $hold(negedge G, posedge D, 1.0, notifier);

    // mpw G-hl NS-hl ()
    $width(negedge G, 1.0, 0, notifier);

    // mpw G-lh NS-lh ()
    $width(posedge G, 1.0, 0, notifier);

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LALM16N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 07:13:57 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LALM1N(D, G, Q, QB);
  input D, G;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc D --> Q
    (D => Q) = (1.0, 1.0);

    // arc D --> QB
    (D => QB) = (1.0, 1.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (1.0, 1.0);

    // arc G --> QB
    (posedge G => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl G-hl ()
    $setup(negedge D, negedge G, 1.0, notifier);

    // setup D-lh G-hl ()
    $setup(posedge D, negedge G, 1.0, notifier);

    // hold D-hl G-hl ()
    $hold(negedge G, negedge D, 1.0, notifier);

    // hold D-lh G-hl ()
    $hold(negedge G, posedge D, 1.0, notifier);

    // mpw G-hl NS-hl ()
    $width(negedge G, 1.0, 0, notifier);

    // mpw G-lh NS-lh ()
    $width(posedge G, 1.0, 0, notifier);

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LALM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 21:11:32 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LALM2N(D, G, Q, QB);
  input D, G;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc D --> Q
    (D => Q) = (1.0, 1.0);

    // arc D --> QB
    (D => QB) = (1.0, 1.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (1.0, 1.0);

    // arc G --> QB
    (posedge G => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl G-hl ()
    $setup(negedge D, negedge G, 1.0, notifier);

    // setup D-lh G-hl ()
    $setup(posedge D, negedge G, 1.0, notifier);

    // hold D-hl G-hl ()
    $hold(negedge G, negedge D, 1.0, notifier);

    // hold D-lh G-hl ()
    $hold(negedge G, posedge D, 1.0, notifier);

    // mpw G-hl NS-hl ()
    $width(negedge G, 1.0, 0, notifier);

    // mpw G-lh NS-lh ()
    $width(posedge G, 1.0, 0, notifier);

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LALM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 07:18:33 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LALM3N(D, G, Q, QB);
  input D, G;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc D --> Q
    (D => Q) = (1.0, 1.0);

    // arc D --> QB
    (D => QB) = (1.0, 1.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (1.0, 1.0);

    // arc G --> QB
    (posedge G => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl G-hl ()
    $setup(negedge D, negedge G, 1.0, notifier);

    // setup D-lh G-hl ()
    $setup(posedge D, negedge G, 1.0, notifier);

    // hold D-hl G-hl ()
    $hold(negedge G, negedge D, 1.0, notifier);

    // hold D-lh G-hl ()
    $hold(negedge G, posedge D, 1.0, notifier);

    // mpw G-hl NS-hl ()
    $width(negedge G, 1.0, 0, notifier);

    // mpw G-lh NS-lh ()
    $width(posedge G, 1.0, 0, notifier);

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LALM3N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 21:17:06 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LALM4N(D, G, Q, QB);
  input D, G;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc D --> Q
    (D => Q) = (1.0, 1.0);

    // arc D --> QB
    (D => QB) = (1.0, 1.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (1.0, 1.0);

    // arc G --> QB
    (posedge G => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl G-hl ()
    $setup(negedge D, negedge G, 1.0, notifier);

    // setup D-lh G-hl ()
    $setup(posedge D, negedge G, 1.0, notifier);

    // hold D-hl G-hl ()
    $hold(negedge G, negedge D, 1.0, notifier);

    // hold D-lh G-hl ()
    $hold(negedge G, posedge D, 1.0, notifier);

    // mpw G-hl NS-hl ()
    $width(negedge G, 1.0, 0, notifier);

    // mpw G-lh NS-lh ()
    $width(posedge G, 1.0, 0, notifier);

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LALM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 07:16:15 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LALM6N(D, G, Q, QB);
  input D, G;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc D --> Q
    (D => Q) = (1.0, 1.0);

    // arc D --> QB
    (D => QB) = (1.0, 1.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (1.0, 1.0);

    // arc G --> QB
    (posedge G => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl G-hl ()
    $setup(negedge D, negedge G, 1.0, notifier);

    // setup D-lh G-hl ()
    $setup(posedge D, negedge G, 1.0, notifier);

    // hold D-hl G-hl ()
    $hold(negedge G, negedge D, 1.0, notifier);

    // hold D-lh G-hl ()
    $hold(negedge G, posedge D, 1.0, notifier);

    // mpw G-hl NS-hl ()
    $width(negedge G, 1.0, 0, notifier);

    // mpw G-lh NS-lh ()
    $width(posedge G, 1.0, 0, notifier);

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LALM6N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 21:11:26 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LALM8N(D, G, Q, QB);
  input D, G;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1), .preset(1'b1),
        .notifier(notifier));

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc D --> Q
    (D => Q) = (1.0, 1.0);

    // arc D --> QB
    (D => QB) = (1.0, 1.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (1.0, 1.0);

    // arc G --> QB
    (posedge G => ( QB +: D )) = (1.0, 1.0);



    // setup D-hl G-hl ()
    $setup(negedge D, negedge G, 1.0, notifier);

    // setup D-lh G-hl ()
    $setup(posedge D, negedge G, 1.0, notifier);

    // hold D-hl G-hl ()
    $hold(negedge G, negedge D, 1.0, notifier);

    // hold D-lh G-hl ()
    $hold(negedge G, posedge D, 1.0, notifier);

    // mpw G-hl NS-hl ()
    $width(negedge G, 1.0, 0, notifier);

    // mpw G-lh NS-lh ()
    $width(posedge G, 1.0, 0, notifier);

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LALM8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 21:16:44 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LEVUDM12N(A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // LEVUDM12N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 07:14:28 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LEVUDM16N(A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // LEVUDM16N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 07:17:38 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LEVUDM1N(A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // LEVUDM1N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 07:13:54 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LEVUDM2N(A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // LEVUDM2N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 07:16:16 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LEVUDM3N(A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // LEVUDM3N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 07:18:34 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LEVUDM4N(A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // LEVUDM4N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 21:17:09 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LEVUDM6N(A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // LEVUDM6N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 21:16:38 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LEVUDM8N(A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (1.0, 1.0);



  endspecify

  `endif // functional //
endmodule     // LEVUDM8N //
`endcelldefine

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:01:38 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive AD42M1N_UDP5(CO, A, B, C, D, ICI);
output CO;
input A, B, C, D, ICI;
table
// A  B  C  D  ICI : CO
   ?  ?  ?  1    1  :  1;
   0  1  0  ?    1  :  1;
   0  0  1  ?    1  :  1;
   1  0  0  ?    1  :  1;
   1  1  1  1    ?  :  1;
   1  1  1  ?    1  :  1;
   1  0  0  1    ?  :  1;
   0  1  0  1    ?  :  1;
   0  0  1  1    ?  :  1;
   0  1  1  0    ?  :  0;
   0  0  0  0    ?  :  0;
   0  0  0  ?    0  :  0;
   1  0  1  ?    0  :  0;
   1  1  0  ?    0  :  0;
   ?  ?  ?  0    0  :  0;
   0  1  1  ?    0  :  0;
   1  1  0  0    ?  :  0;
   1  0  1  0    ?  :  0;
   
endtable
endprimitive



primitive AD42M1N_UDP6(ICO, A, B, C);
output ICO;
input A, B, C;
table
// A  B  C : ICO
   1  ?  1  : 1;
   1  1  ?  : 1;
   ?  1  1  : 1;
   0  0  ?  : 0;
   0  ?  0  : 0;
   ?  0  0  : 0;
   
endtable
endprimitive



primitive AD42M1N_UDP7(S, A, B, C, D, ICI);
output S;
input A, B, C, D, ICI;
table
// A  B  C  D  ICI : S
   0  0  0  0    1  :  1;
   0  0  1  1    1  :  1;
   1  1  1  1    1  :  1;
   0  0  0  1    0  :  1;
   0  0  1  0    0  :  1;
   1  0  0  1    1  :  1;
   1  0  1  1    0  :  1;
   1  0  1  0    1  :  1;
   1  1  0  0    1  :  1;
   0  1  1  0    1  :  1;
   1  1  0  1    0  :  1;
   0  1  0  1    1  :  1;
   1  0  0  0    0  :  1;
   1  1  1  0    0  :  1;
   0  1  1  1    0  :  1;
   0  1  0  0    0  :  1;
   1  0  1  1    1  :  0;
   1  0  1  0    0  :  0;
   0  0  1  1    0  :  0;
   1  1  0  1    1  :  0;
   0  1  1  1    1  :  0;
   0  1  1  0    0  :  0;
   1  0  0  0    1  :  0;
   1  0  0  1    0  :  0;
   1  1  1  1    0  :  0;
   0  1  0  0    1  :  0;
   0  1  0  1    0  :  0;
   1  1  0  0    0  :  0;
   0  0  1  0    1  :  0;
   0  0  0  1    1  :  0;
   0  0  0  0    0  :  0;
   1  1  1  0    1  :  0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:03:37 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive ADCSCM2N_UDP4(CO0, A, B, NCI0);
output CO0;
input A, B, NCI0;
table
// A  B  NCI0 : CO0
   ?  1     0  :   1;
   1  1     ?  :   1;
   1  ?     0  :   1;
   0  0     ?  :   0;
   0  ?     1  :   0;
   ?  0     1  :   0;
   
endtable
endprimitive



primitive ADCSCM2N_UDP5(CO1, A, B, NCI1);
output CO1;
input A, B, NCI1;
table
// A  B  NCI1 : CO1
   ?  1     0  :   1;
   1  1     ?  :   1;
   1  ?     0  :   1;
   0  0     ?  :   0;
   0  ?     1  :   0;
   ?  0     1  :   0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:01:28 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive ADCSOM2N_UDP4(CO0B, A, B, CI0);
output CO0B;
input A, B, CI0;
table
// A  B  CI0 : CO0B
   0  0    ?  :  1;
   0  ?    0  :  1;
   ?  0    0  :  1;
   1  ?    1  :  0;
   1  1    ?  :  0;
   ?  1    1  :  0;
   
endtable
endprimitive



primitive ADCSOM2N_UDP5(CO1B, A, B, CI1);
output CO1B;
input A, B, CI1;
table
// A  B  CI1 : CO1B
   0  0    ?  :  1;
   0  ?    0  :  1;
   ?  0    0  :  1;
   1  ?    1  :  0;
   1  1    ?  :  0;
   ?  1    1  :  0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:06:36 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive ADFCGCM2N_UDP3(CO, A, B, NCI);
output CO;
input A, B, NCI;
table
// A  B  NCI : CO
   ?  1    0  :  1;
   1  1    ?  :  1;
   1  ?    0  :  1;
   0  0    ?  :  0;
   0  ?    1  :  0;
   ?  0    1  :  0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:06:09 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive ADFCGOM2N_UDP3(COB, A, B, CI);
output COB;
input A, B, CI;
table
// A  B  CI : COB
   0  0   ?  : 1;
   0  ?   0  : 1;
   ?  0   0  : 1;
   1  ?   1  : 0;
   1  1   ?  : 0;
   ?  1   1  : 0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:03:58 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive ADFCM2N_UDP3(CO, A, B, NCI);
output CO;
input A, B, NCI;
table
// A  B  NCI : CO
   ?  1    0  :  1;
   1  1    ?  :  1;
   1  ?    0  :  1;
   0  0    ?  :  0;
   0  ?    1  :  0;
   ?  0    1  :  0;
   
endtable
endprimitive



primitive ADFCM2N_UDP4(S, A, B, NCI);
output S;
input A, B, NCI;
table
// A  B  NCI : S
   0  0    0  :  1;
   1  0    1  :  1;
   1  1    0  :  1;
   0  1    1  :  1;
   1  1    1  :  0;
   0  1    0  :  0;
   1  0    0  :  0;
   0  0    1  :  0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:08:10 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive ADFCSCM2N_UDP5(CO0, A, B, NCI0);
output CO0;
input A, B, NCI0;
table
// A  B  NCI0 : CO0
   ?  1     0  :   1;
   1  1     ?  :   1;
   1  ?     0  :   1;
   0  0     ?  :   0;
   0  ?     1  :   0;
   ?  0     1  :   0;
   
endtable
endprimitive



primitive ADFCSCM2N_UDP6(CO1, A, B, NCI1);
output CO1;
input A, B, NCI1;
table
// A  B  NCI1 : CO1
   ?  1     0  :   1;
   1  1     ?  :   1;
   1  ?     0  :   1;
   0  0     ?  :   0;
   0  ?     1  :   0;
   ?  0     1  :   0;
   
endtable
endprimitive



primitive ADFCSCM2N_UDP7(S, A, B, CS, NCI0, NCI1);
output S;
input A, B, CS, NCI0, NCI1;
table
// A  B  CS  NCI0  NCI1 : S
   1  1   1     ?     0  :   1;
   0  0   1     ?     0  :   1;
   0  0   0     0     ?  :   1;
   1  0   1     ?     1  :   1;
   1  0   0     1     ?  :   1;
   0  1   1     ?     1  :   1;
   0  1   0     1     ?  :   1;
   1  1   0     0     ?  :   1;
   1  1   0     1     ?  :   0;
   1  1   1     ?     1  :   0;
   0  1   0     0     ?  :   0;
   1  0   0     0     ?  :   0;
   0  0   1     ?     1  :   0;
   0  1   1     ?     0  :   0;
   0  0   0     1     ?  :   0;
   1  0   1     ?     0  :   0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:02:57 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive ADFCSOM2N_UDP5(CO0B, A, B, CI0);
output CO0B;
input A, B, CI0;
table
// A  B  CI0 : CO0B
   0  0    ?  :  1;
   0  ?    0  :  1;
   ?  0    0  :  1;
   1  ?    1  :  0;
   1  1    ?  :  0;
   ?  1    1  :  0;
   
endtable
endprimitive



primitive ADFCSOM2N_UDP6(CO1B, A, B, CI1);
output CO1B;
input A, B, CI1;
table
// A  B  CI1 : CO1B
   0  0    ?  :  1;
   0  ?    0  :  1;
   ?  0    0  :  1;
   1  ?    1  :  0;
   1  1    ?  :  0;
   ?  1    1  :  0;
   
endtable
endprimitive



primitive ADFCSOM2N_UDP7(S, A, B, CI0, CI1, CS);
output S;
input A, B, CI0, CI1, CS;
table
// A  B  CI0  CI1  CS : S
   1  1    1    ?   0  : 1;
   0  1    ?    0   1  : 1;
   0  1    0    ?   0  : 1;
   1  1    ?    1   1  : 1;
   0  0    1    ?   0  : 1;
   0  0    ?    1   1  : 1;
   1  0    ?    0   1  : 1;
   1  0    0    ?   0  : 1;
   0  0    ?    0   1  : 0;
   1  1    ?    0   1  : 0;
   0  0    0    ?   0  : 0;
   0  1    ?    1   1  : 0;
   1  1    0    ?   0  : 0;
   1  0    ?    1   1  : 0;
   0  1    1    ?   0  : 0;
   1  0    1    ?   0  : 0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:05:48 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive ADFM0N_UDP3(CO, A, B, CI);
output CO;
input A, B, CI;
table
// A  B  CI : CO
   1  ?   1  : 1;
   1  1   ?  : 1;
   ?  1   1  : 1;
   0  0   ?  : 0;
   0  ?   0  : 0;
   ?  0   0  : 0;
   
endtable
endprimitive



primitive ADFM0N_UDP4(S, A, B, CI);
output S;
input A, B, CI;
table
// A  B  CI : S
   1  1   1  : 1;
   0  1   0  : 1;
   1  0   0  : 1;
   0  0   1  : 1;
   0  0   0  : 0;
   1  0   1  : 0;
   1  1   0  : 0;
   0  1   1  : 0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:08:36 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive ADFOM2N_UDP3(COB, A, B, CI);
output COB;
input A, B, CI;
table
// A  B  CI : COB
   0  0   ?  : 1;
   0  ?   0  : 1;
   ?  0   0  : 1;
   1  ?   1  : 0;
   1  1   ?  : 0;
   ?  1   1  : 0;
   
endtable
endprimitive



primitive ADFOM2N_UDP4(S, A, B, CI);
output S;
input A, B, CI;
table
// A  B  CI : S
   1  1   1  : 1;
   0  1   0  : 1;
   1  0   0  : 1;
   0  0   1  : 1;
   0  0   0  : 0;
   1  0   1  : 0;
   1  1   0  : 0;
   0  1   1  : 0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:06:17 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive AN3M0N_UDP3(Z, A, B, C);
output Z;
input A, B, C;
table
// A  B  C : Z
   1  1  1  : 1;
   ?  0  ?  : 0;
   0  ?  ?  : 0;
   ?  ?  0  : 0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:01:33 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive AN4M0N_UDP4(Z, A, B, C, D);
output Z;
input A, B, C, D;
table
// A  B  C  D : Z
   1  1  1  1  : 1;
   ?  ?  ?  0  : 0;
   ?  ?  0  ?  : 0;
   ?  0  ?  ?  : 0;
   0  ?  ?  ?  : 0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:03:21 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive AO22B10M0N_UDP4(Z, A1, B1, B2, NA2);
output Z;
input A1, B1, B2, NA2;
table
// A1  B1  B2  NA2 : Z
    1   ?   ?    0  :  1;
    ?   1   1    ?  :  1;
    ?   ?   0    1  :  0;
    0   0   ?    ?  :  0;
    0   ?   0    ?  :  0;
    ?   0   ?    1  :  0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:02:03 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive AO22B11M0N_UDP4(Z, A1, B1, NA2, NB2);
output Z;
input A1, B1, NA2, NB2;
table
// A1  B1  NA2  NB2 : Z
    1   ?    0    ?  :  1;
    ?   1    ?    0  :  1;
    ?   ?    1    1  :  0;
    0   0    ?    ?  :  0;
    0   ?    ?    1  :  0;
    ?   0    1    ?  :  0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:09:26 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive AO22M0N_UDP4(Z, A1, A2, B1, B2);
output Z;
input A1, A2, B1, B2;
table
// A1  A2  B1  B2 : Z
    ?   ?   1   1  : 1;
    1   1   ?   ?  : 1;
    0   ?   0   ?  : 0;
    ?   0   0   ?  : 0;
    ?   0   ?   0  : 0;
    0   ?   ?   0  : 0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:08:09 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive AOI211M0N_UDP4(Z, A1, A2, B, C);
output Z;
input A1, A2, B, C;
table
// A1  A2  B  C : Z
    ?   0  0  0  : 1;
    0   ?  0  0  : 1;
    1   1  ?  ?  : 0;
    ?   ?  ?  1  : 0;
    ?   ?  1  ?  : 0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:07:46 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive AOI221M0N_UDP5(Z, A1, A2, B1, B2, C);
output Z;
input A1, A2, B1, B2, C;
table
// A1  A2  B1  B2  C : Z
    ?   0   ?   0  0  : 1;
    ?   0   0   ?  0  : 1;
    0   ?   0   ?  0  : 1;
    0   ?   ?   0  0  : 1;
    ?   ?   ?   ?  1  : 0;
    ?   ?   1   1  ?  : 0;
    1   1   ?   ?  ?  : 0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:03:25 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive AOI222M0N_UDP6(Z, A1, A2, B1, B2, C1, C2);
output Z;
input A1, A2, B1, B2, C1, C2;
table
// A1  A2  B1  B2  C1  C2 : Z
    ?   0   ?   0   0   ?  : 1;
    0   ?   0   ?   ?   0  : 1;
    0   ?   0   ?   0   ?  : 1;
    ?   0   0   ?   0   ?  : 1;
    0   ?   ?   0   ?   0  : 1;
    0   ?   ?   0   0   ?  : 1;
    ?   0   0   ?   ?   0  : 1;
    ?   0   ?   0   ?   0  : 1;
    ?   ?   1   1   ?   ?  : 0;
    ?   ?   ?   ?   1   1  : 0;
    1   1   ?   ?   ?   ?  : 0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:09:45 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive BEMXBM2N_UDP5(PB, M0, M1, OA1, OA2, Z);
output PB;
input M0, M1, OA1, OA2, Z;
table
// M0  M1  OA1  OA2  Z : PB
    ?   1    1    ?  0  : 1;
    1   ?    1    ?  1  : 1;
    0   ?    ?    1  1  : 1;
    ?   0    ?    1  0  : 1;
    ?   1    0    ?  0  : 0;
    ?   0    ?    0  0  : 0;
    1   ?    0    ?  1  : 0;
    0   ?    ?    0  1  : 0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:05:01 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive BEMXM2N_UDP5(P, M0, M1, OA1, OA2, Z);
output P;
input M0, M1, OA1, OA2, Z;
table
// M0  M1  OA1  OA2  Z : P
    ?   1    0    ?  0  : 1;
    ?   0    ?    0  0  : 1;
    1   ?    0    ?  1  : 1;
    0   ?    ?    0  1  : 1;
    ?   1    1    ?  0  : 0;
    1   ?    1    ?  1  : 0;
    0   ?    ?    1  1  : 0;
    ?   0    ?    1  0  : 0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:05:16 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive DFEZRM0N_UDP__OUT__(__OUT__, D, E, IQ, RB);
output __OUT__;
input D, E, IQ, RB;
table
// D  E  IQ  RB : __OUT__
   ?  0   1   1  : 1;
   1  1   ?   1  : 1;
   0  1   ?   ?  : 0;
   ?  0   0   ?  : 0;
   ?  ?   ?   0  : 0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:11:41 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive HSDFEQM1N_UDP__OUT__(__OUT__, D, E, IQ, SD, SE);
output __OUT__;
input D, E, IQ, SD, SE;
table
// D  E  IQ  SD  SE : __OUT__
   ?  ?   ?   1   1  : 1;
   ?  0   1   ?   0  : 1;
   1  1   ?   ?   0  : 1;
   0  1   ?   ?   0  : 0;
   ?  ?   ?   0   1  : 0;
   ?  0   0   ?   0  : 0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:17:51 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive MUX3M0N_UDP5(Z, A, B, C, S0, S1);
output Z;
input A, B, C, S0, S1;
table
// A  B  C  S0  S1 : Z
   ?  1  ?   1   0  : 1;
   ?  ?  1   ?   1  : 1;
   1  ?  ?   0   0  : 1;
   ?  ?  0   ?   1  : 0;
   0  ?  ?   0   0  : 0;
   ?  0  ?   1   0  : 0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:17:07 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive MUX4M0N_UDP6(Z, A, B, C, D, S0, S1);
output Z;
input A, B, C, D, S0, S1;
table
// A  B  C  D  S0  S1 : Z
   ?  ?  ?  1   1   1  : 1;
   ?  1  ?  ?   1   0  : 1;
   ?  ?  1  ?   0   1  : 1;
   1  ?  ?  ?   0   0  : 1;
   ?  0  ?  ?   1   0  : 0;
   0  ?  ?  ?   0   0  : 0;
   ?  ?  ?  0   1   1  : 0;
   ?  ?  0  ?   0   1  : 0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:12:48 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive MXB3M0N_UDP5(Z, A, B, C, S0, S1);
output Z;
input A, B, C, S0, S1;
table
// A  B  C  S0  S1 : Z
   ?  ?  0   ?   1  : 1;
   0  ?  ?   0   0  : 1;
   ?  0  ?   1   0  : 1;
   ?  1  ?   1   0  : 0;
   ?  ?  1   ?   1  : 0;
   1  ?  ?   0   0  : 0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:13:59 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive MXB4M0N_UDP6(Z, A, B, C, D, S0, S1);
output Z;
input A, B, C, D, S0, S1;
table
// A  B  C  D  S0  S1 : Z
   ?  0  ?  ?   1   0  : 1;
   0  ?  ?  ?   0   0  : 1;
   ?  ?  ?  0   1   1  : 1;
   ?  ?  0  ?   0   1  : 1;
   ?  ?  ?  1   1   1  : 0;
   ?  1  ?  ?   1   0  : 0;
   ?  ?  1  ?   0   1  : 0;
   1  ?  ?  ?   0   0  : 0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:17:37 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive ND3B1M0N_UDP3(Z, B, C, NA);
output Z;
input B, C, NA;
table
// B  C  NA : Z
   ?  0   ?  : 1;
   0  ?   ?  : 1;
   ?  ?   1  : 1;
   1  1   0  : 0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:20:05 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive ND3M0N_UDP3(Z, A, B, C);
output Z;
input A, B, C;
table
// A  B  C : Z
   ?  0  ?  : 1;
   0  ?  ?  : 1;
   ?  ?  0  : 1;
   1  1  1  : 0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:13:13 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive ND4B1M0N_UDP4(Z, B, C, D, NA);
output Z;
input B, C, D, NA;
table
// B  C  D  NA : Z
   ?  ?  ?   1  : 1;
   ?  ?  0   ?  : 1;
   ?  0  ?   ?  : 1;
   0  ?  ?   ?  : 1;
   1  1  1   0  : 0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:19:32 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive ND4B2M0N_UDP4(Z, C, D, NA, NB);
output Z;
input C, D, NA, NB;
table
// C  D  NA  NB : Z
   ?  ?   ?   1  : 1;
   ?  0   ?   ?  : 1;
   ?  ?   1   ?  : 1;
   0  ?   ?   ?  : 1;
   1  1   0   0  : 0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:18:07 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive ND4M0N_UDP4(Z, A, B, C, D);
output Z;
input A, B, C, D;
table
// A  B  C  D : Z
   ?  ?  ?  0  : 1;
   ?  ?  0  ?  : 1;
   ?  0  ?  ?  : 1;
   0  ?  ?  ?  : 1;
   1  1  1  1  : 0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:18:44 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive NR3B1M0N_UDP3(Z, B, C, NA);
output Z;
input B, C, NA;
table
// B  C  NA : Z
   0  0   1  : 1;
   ?  1   ?  : 0;
   1  ?   ?  : 0;
   ?  ?   0  : 0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:16:18 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive NR3M0N_UDP3(Z, A, B, C);
output Z;
input A, B, C;
table
// A  B  C : Z
   0  0  0  : 1;
   ?  1  ?  : 0;
   1  ?  ?  : 0;
   ?  ?  1  : 0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:16:05 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive NR4B1M0N_UDP4(Z, B, C, D, NA);
output Z;
input B, C, D, NA;
table
// B  C  D  NA : Z
   0  0  0   1  : 1;
   ?  ?  ?   0  : 0;
   1  ?  ?   ?  : 0;
   ?  1  ?   ?  : 0;
   ?  ?  1   ?  : 0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:13:44 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive NR4B2M0N_UDP4(Z, C, D, NA, NB);
output Z;
input C, D, NA, NB;
table
// C  D  NA  NB : Z
   0  0   1   1  : 1;
   ?  ?   ?   0  : 0;
   1  ?   ?   ?  : 0;
   ?  ?   0   ?  : 0;
   ?  1   ?   ?  : 0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:13:45 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive NR4M0N_UDP4(Z, A, B, C, D);
output Z;
input A, B, C, D;
table
// A  B  C  D : Z
   0  0  0  0  : 1;
   ?  ?  ?  1  : 0;
   ?  1  ?  ?  : 0;
   ?  ?  1  ?  : 0;
   1  ?  ?  ?  : 0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:16:20 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive OAI221M0N_UDP5(Z, A1, A2, B1, B2, C);
output Z;
input A1, A2, B1, B2, C;
table
// A1  A2  B1  B2  C : Z
    ?   ?   ?   ?  0  : 1;
    ?   ?   0   0  ?  : 1;
    0   0   ?   ?  ?  : 1;
    ?   1   1   ?  1  : 0;
    ?   1   ?   1  1  : 0;
    1   ?   ?   1  1  : 0;
    1   ?   1   ?  1  : 0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:14:30 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive OAI222M0N_UDP6(Z, A1, A2, B1, B2, C1, C2);
output Z;
input A1, A2, B1, B2, C1, C2;
table
// A1  A2  B1  B2  C1  C2 : Z
    ?   ?   ?   ?   0   0  : 1;
    0   0   ?   ?   ?   ?  : 1;
    ?   ?   0   0   ?   ?  : 1;
    1   ?   1   ?   1   ?  : 0;
    1   ?   ?   1   ?   1  : 0;
    ?   1   1   ?   ?   1  : 0;
    1   ?   ?   1   1   ?  : 0;
    1   ?   1   ?   ?   1  : 0;
    ?   1   ?   1   1   ?  : 0;
    ?   1   ?   1   ?   1  : 0;
    ?   1   1   ?   1   ?  : 0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:14:09 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive OAI22B10M0N_UDP4(Z, A1, B1, B2, NA2);
output Z;
input A1, B1, B2, NA2;
table
// A1  B1  B2  NA2 : Z
    ?   0   0    ?  :  1;
    0   ?   ?    1  :  1;
    1   1   ?    ?  :  0;
    ?   1   ?    0  :  0;
    1   ?   1    ?  :  0;
    ?   ?   1    0  :  0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:14:19 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive OAI22B20M0N_UDP4(Z, B1, B2, NA1, NA2);
output Z;
input B1, B2, NA1, NA2;
table
// B1  B2  NA1  NA2 : Z
    ?   ?    1    1  :  1;
    0   0    ?    ?  :  1;
    ?   1    0    ?  :  0;
    1   ?    ?    0  :  0;
    1   ?    0    ?  :  0;
    ?   1    ?    0  :  0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:21:37 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive OAI22M0N_UDP4(Z, A1, A2, B1, B2);
output Z;
input A1, A2, B1, B2;
table
// A1  A2  B1  B2 : Z
    0   0   ?   ?  : 1;
    ?   ?   0   0  : 1;
    ?   1   ?   1  : 0;
    1   ?   ?   1  : 0;
    1   ?   1   ?  : 0;
    ?   1   1   ?  : 0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:19:12 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive OAI31M0N_UDP4(Z, A1, A2, A3, B);
output Z;
input A1, A2, A3, B;
table
// A1  A2  A3  B : Z
    ?   ?   ?  0  : 1;
    0   0   0  ?  : 1;
    ?   ?   1  1  : 0;
    1   ?   ?  1  : 0;
    ?   1   ?  1  : 0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:19:24 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive OAI32M0N_UDP5(Z, A1, A2, A3, B1, B2);
output Z;
input A1, A2, A3, B1, B2;
table
// A1  A2  A3  B1  B2 : Z
    ?   ?   ?   0   0  : 1;
    0   0   0   ?   ?  : 1;
    1   ?   ?   ?   1  : 0;
    ?   ?   1   1   ?  : 0;
    1   ?   ?   1   ?  : 0;
    ?   1   ?   1   ?  : 0;
    ?   1   ?   ?   1  : 0;
    ?   ?   1   ?   1  : 0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:19:54 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive OAI33M0N_UDP6(Z, A1, A2, A3, B1, B2, B3);
output Z;
input A1, A2, A3, B1, B2, B3;
table
// A1  A2  A3  B1  B2  B3 : Z
    0   0   0   ?   ?   ?  : 1;
    ?   ?   ?   0   0   0  : 1;
    ?   ?   1   1   ?   ?  : 0;
    ?   ?   1   ?   ?   1  : 0;
    1   ?   ?   ?   ?   1  : 0;
    1   ?   ?   1   ?   ?  : 0;
    1   ?   ?   ?   1   ?  : 0;
    ?   1   ?   1   ?   ?  : 0;
    ?   1   ?   ?   ?   1  : 0;
    ?   1   ?   ?   1   ?  : 0;
    ?   ?   1   ?   1   ?  : 0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:15:13 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive SDFEM0N_UDP__OUT__(__OUT__, D, E, IQ, SD, SE);
output __OUT__;
input D, E, IQ, SD, SE;
table
// D  E  IQ  SD  SE : __OUT__
   ?  ?   ?   1   1  : 1;
   ?  0   1   ?   0  : 1;
   1  1   ?   ?   0  : 1;
   0  1   ?   ?   0  : 0;
   ?  ?   ?   0   1  : 0;
   ?  0   0   ?   0  : 0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:14:38 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive SDFEQBM0N_UDP__OUT__(__OUT__, D, E, IQ, SD, SE);
output __OUT__;
input D, E, IQ, SD, SE;
table
// D  E  IQ  SD  SE : __OUT__
   ?  ?   ?   1   1  : 1;
   ?  0   1   ?   0  : 1;
   1  1   ?   ?   0  : 1;
   0  1   ?   ?   0  : 0;
   ?  ?   ?   0   1  : 0;
   ?  0   0   ?   0  : 0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 19:15:31 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive SDFEZRM0N_UDP__OUT__(__OUT__, D, E, IQ, RB, SD, SE);
output __OUT__;
input D, E, IQ, RB, SD, SE;
table
// D  E  IQ  RB  SD  SE : __OUT__
   1  1   ?   1   ?   0  : 1;
   ?  ?   ?   ?   1   1  : 1;
   ?  0   1   1   ?   0  : 1;
   ?  ?   ?   0   ?   0  : 0;
   ?  0   0   ?   ?   0  : 0;
   0  1   ?   ?   ?   0  : 0;
   ?  ?   ?   ?   0   1  : 0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:19:53 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive XNR3M0N_UDP3(Z, A, B, C);
output Z;
input A, B, C;
table
// A  B  C : Z
   0  0  0  : 1;
   1  0  1  : 1;
   1  1  0  : 1;
   0  1  1  : 1;
   1  1  1  : 0;
   0  1  0  : 0;
   1  0  0  : 0;
   0  0  1  : 0;
   
endtable
endprimitive

/*****************************************************************************/
/*                                                                           */
/*  SiliconSmart CR 2005.05, build 15 production                             */
/*  Created:  Wed Aug  3 05:20:40 2005 by weiluen                            */
/*    for Verilog Simulator:  verilog-xl                                     */
/*                                                                           */
/*****************************************************************************/

`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive XOR3M0N_UDP3(Z, A, B, C);
output Z;
input A, B, C;
table
// A  B  C : Z
   1  1  1  : 1;
   0  1  0  : 1;
   1  0  0  : 1;
   0  0  1  : 1;
   0  0  0  : 0;
   1  0  1  : 0;
   1  1  0  : 0;
   0  1  1  : 0;
   
endtable
endprimitive

// CR default primitives
// All cells assume preset and clear are active low


///////////////////////////////////////////////////////////////////////////
// This dff cell has a reset priority over preset

primitive udp_dff_p0(q, d, clk, clear, preset, notifier);
	output q;
	input  clk, clear, d, preset, notifier;
	reg q; /* declaring output as reg*/
	
	table
	// d  clk  clear  preset  notifier : state : q
           0   r    ?      1     ?    : ?  :  0  ; // clock in 0
           1   r    1      ?     ?    : ?  :  1  ; // clock in 1

           1   *    1      ?     ?    : 1  :  1  ; // reduce pessimism
           0   *    ?      1     ?    : 0  :  0  ; // reduce pessimism

           ?   f    ?      ?     ?    : ?  :  -  ; // no changes on negedge clk
           *   b    ?      ?     ?    : ?  :  -  ; // no changes when in switches

           ?   ?    0      ?     ?    : ?  :  0  ; // reset output; dominate

           ?   b    1      *     ?    : 1  :  1  ; // cover all transistions on set_
           1   x    1      *     ?    : 1  :  1  ; // cover all transistions on set_

           ?   ?    1      0     ?    : ?  :  1  ; // set output

           ?   b    *      1     ?    : 0  :  0  ; // cover all transistions on clr_
           0   x    *      1     ?    : 0  :  0  ; // cover all transistions on clr_

`ifdef SMC_NFORCE	
	   ?   ?     ?      ?        *     :   ?   : x ;  // on any notifier event output x
`else
	   ?   ?     ?      ?        *     :   ?   : - ;  // ignore notifier changes in functional mode
`endif
	endtable
endprimitive

module dff_p0(q, d, clk, clear, preset, notifier);
   output q;
   input  clk, clear, d, preset, notifier;

   udp_dff_p0 D1(q, d, clk, clear, preset, notifier);
endmodule // dff_p0

///////////////////////////////////////////////////////////////////////////
// This cell has a preset priority over reset

primitive udp_dff_p1(q, d, clk, clear, preset, notifier);
	output q;
	input  clk, clear, d, preset, notifier;
	reg q; /* declaring output as reg*/
	
	table
	// d  clk  clear  preset  notifier : state : q
           0   r    ?      1     ?    : ?  :  0  ; // clock in 0
           1   r    1      ?     ?    : ?  :  1  ; // clock in 1

           1   *    1      ?     ?    : 1  :  1  ; // reduce pessimism
           0   *    ?      1     ?    : 0  :  0  ; // reduce pessimism

           ?   f    ?      ?     ?    : ?  :  -  ; // no changes on negedge clk
           *   b    ?      ?     ?    : ?  :  -  ; // no changes when in switches

           ?   ?    ?      0     ?    : ?  :  1  ; // set output; dominate

           ?   b    1      *     ?    : 1  :  1  ; // cover all transistions on set_
           1   x    1      *     ?    : 1  :  1  ; // cover all transistions on set_

           ?   ?    0      1     ?    : ?  :  0  ; // reset output

           ?   b    *      1     ?    : 0  :  0  ; // cover all transistions on clr_
           0   x    *      1     ?    : 0  :  0  ; // cover all transistions on clr_
`ifdef SMC_NFORCE	
	   ?   ?     ?      ?        *     :   ?   : x ;  // on any notifier event output x
`else
	   ?   ?     ?      ?        *     :   ?   : - ;  // ignore notifier changes in functional mode
`endif
	endtable
endprimitive

module dff_p1(q, d, clk, clear, preset, notifier);
   output q;
   input  clk, clear, d, preset, notifier;

   udp_dff_p1 D1(q, d, clk, clear, preset, notifier);
endmodule // dff_p1



///////////////////////////////////////////////////////////////////////////
//

primitive udp_inv_clr0 (qn, clr, pre, inp);
	output qn;
	input  clr, pre, inp;

	table

	//  	clr 	pre 	inp	: qn
		0	0	?	: 0;
		1	?	0	: 1;
		1	?	1	: 0;
		?	1	0	: 1;
		?	1	1	: 0;
		x	x	1	: 0;
		x	x	0	: 1;
	endtable
endprimitive

module inv_clr0 (qn, clr, pre, inp);
   output qn;
   input  clr, pre, inp; 

   udp_inv_clr0 (qn, clr, pre, inp);
endmodule // inv_clr0


///////////////////////////////////////////////////////////////////////////
//

primitive udp_mux21 (q, data1, data0, dselect);
    output q;
    input data1, data0, dselect;

// FUNCTION :  TWO TO ONE MULTIPLEXER
table
//data1 data0 dselect :   q
        0     0       ?   :   0 ;
        1     1       ?   :   1 ;

        0     ?       1   :   0 ;
        1     ?       1   :   1 ;

        ?     0       0   :   0 ;
        ?     1       0   :   1 ;
endtable
endprimitive


module mux21 (q, data1, data0, dselect);
   output q;
   input  data1, data0, dselect;

   udp_mux21 m1(q, data1, data0, dselect);
endmodule // mux21

///////////////////////////////////////////////////////////////////////////
//

primitive udp_ldlatch_p0(q, d, en, clear, preset, notifier);
	output q;
	input  d, en, clear, preset, notifier;
	reg q;

	table
	// d  en  clear	 preset	 notifier : state : q
           1  1    1     ?        ?       : ?  :  1  ; // 
           0  1    ?     1        ?       : ?  :  0  ; // 
           1  *    1     ?        ?       : 1  :  1  ; // reduce pessimism
           0  *    ?     1        ?       : 0  :  0  ; // reduce pessimism
           *  0    ?     ?        ?       : ?  :  -  ; // no changes when in switches

           ?  ?    0     ?        ?       : ?  :  0  ; // reset output : reset dominate

           ?  0    1     *        ?       : 1  :  1  ; // cover all transistions on set_
           1  ?    1     *        ?       : 1  :  1  ; // cover all transistions on set_

           ?  ?    1     0        ?       : ?  :  1  ; // set output

           ?  0    *     1        ?       : 0  :  0  ; // cover all transistions on clr_
           0  ?    *     1        ?       : 0  :  0  ; // cover all transistions on clr_
`ifdef SMC_NFORCE	
	   ?  ?    ?     ?        *       : ?  :  x ;  // on any notifier event output x
`else
	   ?  ?    ?     ?        *       : ?  :  - ;  // ignore notifier changes in functional mode
`endif
	endtable
endprimitive

module ldlatch_p0(q, d, en, clear, preset, notifier);
   output q;
   input  clear, preset, d, en, notifier;

   udp_ldlatch_p0 P1 (q, d, en, clear, preset, notifier);
endmodule // ldlatch_p0

///////////////////////////////////////////////////////////////////////////
//

primitive udp_ldlatch_p1(q, d, en, clear, preset, notifier);
	output q;
	input  clear, preset, d, en, notifier;
	reg q;

	table
	// d  en  clear	 preset	 notifier : state : q
           1  1   1   ?   ?   : ?  :  1  ; // 
           0  1   ?   1   ?   : ?  :  0  ; // 
           1  *   1   ?   ?   : 1  :  1  ; // reduce pessimism
           0  *   ?   1   ?   : 0  :  0  ; // reduce pessimism
           *  0   ?   ?   ?   : ?  :  -  ; // no changes when in switches
           ?  ?   ?   0   ?   : ?  :  1  ; // set output
           ?  0   1   *   ?   : 1  :  1  ; // cover all transistions on set_
           1  ?   1   *   ?   : 1  :  1  ; // cover all transistions on set_
           ?  ?   0   1   ?   : ?  :  0  ; // reset output
           ?  0   *   1   ?   : 0  :  0  ; // cover all transistions on clr_
           0  ?   *   1   ?   : 0  :  0  ; // cover all transistions on clr_
`ifdef SMC_NFORCE
	   ?   ?    ?      ?        *     :   ?   : x ;  // on any notifier event output x
`else
	   ?   ?    ?      ?        *     :   ?   : - ;  // ignore notifier changes in functional mode
`endif
	endtable
endprimitive

module ldlatch_p1(q, d, en, clear, preset, notifier);
   output q;
   input clear, preset, d, en, notifier;

   udp_ldlatch_p1 P1 (q, d, en, clear, preset, notifier);
endmodule // ldlatch_p1